`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
c4q0gy3SzyhhckDi/m2sCHEg71u5lxr9H1vV9ouGQEGV3nLKmOk5yZIrSjPIoXSSyk9p1ZKLrmkB
TiFTKvcrzg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
REt97Ap4rm2nsvnOnsIRXZD465mWqnJSqP2D9OtzP5PtnVMKQRSg0GJAe51zopUuItBBuYdO+2qB
EaALk55wHxUSfAfyCq7KVoBbeFmzJY7hDHAq3JIslggkKK3qB9PV2SVfj+6Jk8y6uujjQb9iq5bs
fImmvi16ao2mz1pqPJ4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FBenFuPBh0Ptgf14Ex1U5CcRJ23qr6l/dap6TJK+ypHJDHJ1bKrlr6rx7Db/1Crd2ru3yQkv1Neu
7Eiq+yvhZv9VJKQFxPevdsRVIG4dSnY6TiGjhDMQrT8g9F5+WuKC/h6T9lMJFQ02ctmhbxRX6CWg
o5WJVVgfaqQRVDZiyfZxggLQ9qTK+OPqL4q46t+peV2bZrFQXjQbAOTTGm4trKKpffZQUgmx793q
ehDW5vCIuJroonxsmOofmV5GSpao4COmqvjNf6bpQHKow9TkLhn9XG68Iz1cCOXYKUI80pB/5WAq
THRG13MBHkE24/tDaavBdcV8T7UGkYaYs1/Y/Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xUTFAuNDBAX7+LLAcpbupN25K1dkz24OrtZPhDjPOe52lqY88up1J0en+rAyCofVbDif5SmPype7
aXr3CDqS0yCfEtgkIdszMu5TqiDFo5QRVdQJaqNKhRf8UF3njPx4uifpcpJ1OmwfqQ+FDo1S2qFD
h/VGBSGm/mJy8i3KQIk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kSf866Twzle8aoPcriukhSamNwggln16bvz77fjv6GgvYfzg+2WofrMbcCi0Uy8EOhM/+cNIh1cB
R7V6y2vIPvzFiYv/GiG85ufyY/fP0GFRpOUsfsQyWtFI6zdJ7Wh88R/bx9SaRZZqMF53cLSz1J1R
m1mYzqAVakWgO+p3+JKcpm5Ef0tXCLqNxY87xQE9km5RkZYQwRtUCTt02KeJ5ktmJXKL60MVGFWc
4/4Z2GpL56d9kKWhIZ7DQR8nSGvkOv97IYmFOAEFtZzcKX5EEfnTvNghSNm7e/rbFdUK6LedIt5G
PlzlrPY9MrmM8Ehnq0trQ+t+7Xh1l5/LkOzPNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23776)
`protect data_block
3bSOmz+xdKOeL2nMpt0bVkLHQP7S68ssPxPtobaMqmF7kcY2DubtzCNl77gkkVCHVxEynzxufSpU
OGlHv+YJlykooewOHowP9HahVqiKPiO/I0YB3gaVK6gBGYQUHsfhCUe75FuKb6CeORCqmFuAR+N+
kyv4HnouskU+6lQNabAowUToMSW1/Bl4Bzn/tiogTvsY7j+VoGBLp+UoEV2Q+rpfiH6w2joaIP3n
9OR7XdF9Rno/2upxreuwFO/JlWCcJ2LSI6roGl2bCjI2kbeJXRulHUTQRGlYl4UN5FxmhEm1uc48
SbVxZRStcNiGKCFsjliTYcT7awgCCQKpxFApx//x5YBnUa4jeqdMjKlZAfo0hGQhtCOwzDfSvo3X
kmNeD02H2IpcnDdvcJLzVhvz1VTdjUlNuq6ckCPyDN9zkpJC5coOI/8BW3FDzD0lYOAjDnI0qvIY
dzr3uchfnGS7CaRYETB22YdMuLkLwb7U4A4ZUWKnrtquiH711HV4TrjwFga5mDbgWLvcfYNmErTf
bHeafG+5RMmOHvbt3lu6tEkwvWWhNE/isP1JoYbMkxX8aEijMA4DEvgeJNhwbL4f+8LG1/E5zYOc
ldOsXWaT5f6ML7zzhS7twEf+LUbQmmNMawkEw9JN6KyhDyzXSfTsizQkNBCZyBhvHqTzQr6pI5eR
C9Slhldn9VaV3AlD8mOFFKbTyDtygZtnDLnlwro/2X/AuJ+1JQEpDCupFUMHrZNi51Hk5ensdLKd
V1stys2HKAKfnFwDInpN4XoXq0vuBQ6k1Qs4F711qJ2CGM29uRDs+viucps785+gb4P+3RsVwXJI
r5kZ5V7/BXtGEluNGZsixdYk/WGxHBuJhmmrdWmQOzhG/6RhVDzocxMJiVGdxSgextnm7Y+D1sZf
Xns21SBUv5/eBlORtysQxUMH9zx7G3LrlRkB8kkx2dVzmoRRBp6DhlqgzktzrUTxd+d1O3lxjOr6
4/frjD3bJrN/XsDA0JADvTvB5+n3/qhmR35Hlx9UZocBTLj1l6mfrkz4iLDuAkoCc5EcgYQ2Lbt9
sQsl+c+H1wU/UIEQBxOFkON2uIObkjwWw0rveqIZ/NPaZjtdcw7R2NP/UKRRFENQvpaDLgWy0Qj9
UOx4r1DGYKWMadAVQfidaSYwvECK0zrrG9S3mnJJt+JEeplOqHowq4gJPaMJjvSoiquVbgI/z/WZ
YYqfYont1I6dh2QwGJN0pkLLAswOnm5E8EiODzr7TK73nkPatrSuk3MUonvecjU4ajrcnExv7Yzr
2gH9b9YxEu/HOjQZoGziu3dJb+53hF0Bu99uPntYvLZ52iNiWM8YLIG4Vc8sGdg9ViN84WAunJpE
hJLzO3PdPcmgHYCnauoWE+n0FKGqL+nFHIqQaaAwU84wYl26dcFSn8SpYuYb3yi8y2USBHSAg5DC
TUlz2Ef8jcnHpv+uxpuO02tw2JpUKDn/BGsmc0Slp0gyz1JhvQ8cmfuXgTi7v+ILzS4bUbIKI5ZP
yJKCrjUK9bXSC/kWkp7/K0rXCsg2bNhaAm9A0F3vTc30bwiqqHhONkB5gHyGK09s6erZKhDpL1Fm
yFxhU9uQ4OIhqIS2ek9DwZ5nb5eDx+xI/NZfOC1F0SpNhC/XudTzPezArtOQ8HSQeL6IIOg/83+A
pF0rVPWLis1J3LrHyrIyhWr4B1O1q202ctDuxUYJUyz9eb/rhJbEG7DpiolJKozt4+wCH3sKZXzX
dw+6AUSEnpQ9hVO1ruMLWaK1J8SbRxxrYVj/kna5gk/bEPHgqrq3MvJ/dCgbp5fYkUoTXJCI6yEb
O6RvzHdUm52U3hPqkOcXkKnfGigczIPDWEDU+84UUCJUH0bcvCffVjGwz4jTNlqwlz6YP7qQrCHZ
cWL1tvoGGYejmuZAAB4wfD9aDQ10yKC8EFfVPOA+NsoaBKpePrb5BkUxxY60+ajWOejJkeQQmTNt
scdvpF/FBmYsljRu1Qjk4u8kzjoXAuQU8riohTrnPjvISkKlQoVDqCmuN68TbM+NqSbld+BojzVT
2/ZrV0IoZDrAt8Oj+LMK0TF2rQSKKPm/IMEAyLJf9Pih5EIJ9XAXtm64PggGs311BZO2FwUMa2Cz
T6pSbpr8Hdx4AbKbFS8GqNlzQ7z1Uul52/fv5UjkW6mQmE0RnUdAz0TnDiDCFKXtrzhmtT2w2nWr
uNhfpXIu9vHdmp2rurcldL+OMJLLUSke0bi7s3xXovVXnkHQlCfB+gqyr6ZNv5N7zmhtdVCP7yWz
hqCbAHxABlusm2c1VlS6Jgj7p74iMfVeqLDvemkjrGrYHWTAA2F3tuBQwKNhV/Zahwi9l1Nda+HK
rUCbRQmcL62wMBXaICTn/DMJDSukt+oLg/VHITqmRCNvcln3NAarMtGHWPB1DYBf5QnD8XMHjsQ+
5l0JKJHlyaw8VZ1T50jwYVvhEn5NxlZ0Nyg8oGiEFhh5w/sET7vlRUrwpcYiiOn8PT01tkJmX/+I
zsjONmitx5ez35mzf30HxwZRZl9EvOg0mzVclpXVYQBgqy4pV4w1OtxTez2LxH4SkSgUkexO29wU
ZH43vPNgSwco18Td9Hn7vmypNi2pxe7AQh8G33NmaE4uFhsxNY3/JNsufXasDQZganVciKcNzq7H
obRRXFXvnba6hBGuRnnArFaG6/CX4poCVYXs0a/YrqRm1yi7onq9n4ktGaBNqE+Ie8CT/sZo5SC0
ZcUTMEFMSzu+Guv9ElxWwl2EuL9SYFZMSNT4wlUZLLliZ1pf95SMqWi7s+UIfYfa/NVqLAowX2R+
XYBYxbYUJc1vON8VAINABUtyndox0QjE0/vsBIxc8DK+wsZqXxIaLTZDjh6UXHbpWDJ/EkNhZ1gv
rsJQtw0MFEPN2kd2bnFEpkGIrg/03DDC9ANyIs4YQgGiJ8nXvzTN1YeH95xdiM5Ye94IHmYfOlpe
+SCBIjg7XOYx74OoJ9ftiE2C4POEUTX2y187fD0RiPhlmHpOPxkat1N8nn78auFsjzI5zCW0VJnh
fqWMCYJ4IYJ99b3x0+HsW6Dr9x+UyE1jU+YCBgeshlnCgntyK4doWO647GTJyi6brlUcpTuVIarh
D7Z0xwEeiwgx/lvokXp6TEbM/WTlbKCcLeb/IQFMUJgwH/HdTm1feFFS+QVYzog4sO9Q2Fe5YghH
jiIRqObvkAIFjqfZPijUxarNxSjrqYFS8CYufeyc4Do5zFdq72NSlhMOz4vGghGVfRdRiLnQ68l+
GNb/gqLIMPJGwO6ubDGhFFTmAFjOPmux/0CkJCDRHI6J9js26N3UY5eXfnIW4JvlTI9T97Jy33gN
T6trL/E7UirqtFR7ilh0rDxOqIbT/ZykMHXpNZCES3jZJx2oKgFtYmzHth8oV+lx4DXXtFcvCowy
LCDhbF7zypQlsYo0e9+7ciR4rwVoly4caW8yK83oOOpTeGFiAAperX31If1cYmBBejMJLkTJPhA2
/TqmEZ78jNsshuAZHA9aUw2SK0diAn+zLvSRLmOqzQxq2gB2KWRIeGlJTB//BohR9CiNUzZ88XyV
DuYr8dF3fOwv/9yiROhuVmhxO/lGwCD8va6yy2XVTXwLORCj9m+dmnQF9uZR5FrNndQih6u3/8IF
fwnr7Tqqkta3fIKbOl08Yo37EgTjSqRCxDvT7IXRC4n4iu5MRt0IpIqdQeSZUIgBrvgqz2yzl2Cz
6DNyZWlayTuLJTSgoi0zZgNuNnPJgHnNMpRg5OdcTnULJ9X9FCaPMcObUpx1Z03mOjRtHjEHM3vl
jAu8gSUQwAhzZkdatGLh3Fa65kddZRbquLoTc8XivRchETy71zXVjabsBPc1tDzAyGgaYGLsnj9i
Mh2MOA4ZBD2yIFPNQhJYXwVhpmWroYIzq8SuZXBbVfgK2DGxdAez5rOmQcb5jtVGkbsbROORlkr6
2vUReBjRngDuHNn9DpVPwqkACq4eFHFhVnKX3iJOCB99gCaBmGRaADa9hAbleGOPcLhugbzIZXA9
7R+K8zYzK9J5mKLVi2OeeUE6ckiia3/IHEhDVKxNZacdpelL3W4djWHg5b7FDgMUiRWyMWE89IOM
zcFvVs+sQ6SAVzX4nukoA3hgTRY5Rkivz7ZV9MmL8VfnivGZGZdiIQcAWG2wmRdE7u/n+U0wUYe0
Ua7dqmMoBElYLbIQ2adTvVQvOiYIwlp0vSNjCGrISG7UQsHiA2tPDBF4aQ6l7f+B/OvXOypixjz/
lh5OonudZWdzSCaCeSCH/h7zTQlBVPJcWsaT9cJjk/uHLdqKUOIHNQtbNMSn6xTxgXe4o5UrWcF8
V4Hsfpje4tajvInZryP/ZxkU1Pi/PrPzrEgWwXEfnquRbfzEyh1U0FiIqk9kwsmrpyh74F5LvZGI
I7OMBhSbbPBa29J1DL9fR9bAk0Xx8f9pVVI4GxKNMcPF+c9MJfYCqVrs0qHIIYA18KAwNPB0z1PT
R6u6RqrLmo+9LuvlcLlpgMkKe3mafv5fQCCM0iVdWhQrq+Z0NM+KGdqXuvDMb+qSe8EI6pUoLf5U
JWpStKpaQiDvSG0rINfNjAkg2f4SVuFfsapjVuiZgTIJ0RN0MvE9cEbAawXhp6aWP65YJBbrjmeF
oeqBc2+HWL0ULQJbXpHz4Y4uqPDT6MgrudfzBGvOQ8w3jdRPdgXS4B9pR/8M/bhS1Cv64bVHRFen
807nBxIwFvEvBsvRUwpzReumS7DEIuZbFibCOe0SjQP8/YoVezoQmJrV4TeCk7h8jWqKiLl8tDMR
+d4nHx8CZ4im2vL4Dlm7xvxJtO0/Il8R8kfutujibYTMs6TLIqw2GFf4ajCak+4C9SNhqddkKTPA
iNy/SEf81HpazU6c8a1DT8k7F0GhCBOfwh/tA3PKZYQX5INTd5hEUDG46tUMUTbAFfnMJXChAKyw
lfLDWaLh4YvF8J7NXunP4omKs9vEisOn3KlgZ68smB/BvMg3iasGIY9VXsENtR3IxpY7vMx1oA99
5q7Q9m2oOcTtmLYyh2NSb3TsSH7GT2cPzBe4jRH0W4kOqNFLnW7Kc5KfUn+PKirHIG30cA+u8tBT
NZSMLP+xC5tQ1Jn6CFFhNr1ZwQ8aywL5kv01eRye9JNB4okhZBtKkM7+WcHE2k0vcSy7Z1szlopP
XeoV8BDxd7WnM0P46PKJJddCHsIqAY26NGXFOyr2Kto3ycK+AETNTuGIQWtm1lJpPiVlukmoOkqT
CSUx6gNK/cb2eHKN2aI7oKvqxKOd7x9+I9rxAJmpORAcpH7O7HdAyt4xy8uWumrWhVwAyGnlc6AE
pKQb1cv145+UagzJ/FJh1y/l6e7QZs/moBBmYc7sipybn2GXjjwhItzlwVUiTCwR6Iym1ZHYGQJB
AAlFktnayxFrOAKXzEa0kjKfzYwQZw9cwsQ4XriqIT8fVduOEaohOvndc4A0Nxj7DpMFPMyD+BDY
M+/kw8JUlJ9XRLyr3P9MKZgxq5u0LoEdZIqOIlvIPe9HpQxNPB9FVhQYtRCYXaIcaVJwYetzOLP0
iVt6yN5e5EsyvtNmLY0tU+x4FgyXOp1cT5qkRea75V3Euh38ZW2Sfb14ARRou/qRuBnM/Ea06cxx
s7iivuHv4vP03CNPASCanePw5d25D6tmdo8urQZEezKxuiylcTGzeJxJYTK2tAgZijA1Vgujfl8O
YenqytQVc0PZm5m/1DjlrvD8oHYei040HQIZ7ikDam1CfU45X6+KfI99y+r+7yj93L+I3kAjCBub
y8RRcib5wkpu1i+SQFvH5k9+jFVqIyFOF/Xh2tTJGfWxwTEGKbFrdvZPpFXZiGGQ3NcvhaOYNOF1
dPNpM0eypURYlk5yFQSQgXfPaIxYJB4KIlEAJg92OouZYm3meOktt9AMqBnf7Mf1uP3mgN8JrVfT
EnO+7aAiI9BCMME1o9m2k491p2i+88zwjDKpalx57/L5ENIp3W9IBcyZ2hMPhBycyp04fDbss29l
55IgbAz/1DLNdyETNZCy4TMVvB8k9/0H8E5x1mYHLQwWFFNJ23NFS9LIthKEl5QuJAAqHwZoMIf1
PbrVmh7cDvUATe2rfgYPyycEabc7IcXgyi7hXbFvLhE9w+0qriE21GdCeKJsIsLjnEJshkmYlrmL
jcwQJsacfXxOeNOZkNh6mIt39Z/TvPXp0Q2wtWgWtrdfc8zD9mV8bcq1JJDyZVrmVxvy4fxOcxo/
o0vRF6Ho9SAdf4u4ki4g6xZH0WayaqQQQaRpF85ILloscUpQKvOYTuf/JQcRycxe2sOWx/yfMNHj
gjtkvrhKn9yuQZMFGwEhiuK6dR3ww/f4G/sVNNsw2apJo+lFJR3Rd1oP8OrymiNs/jHAjX3DSPeh
OfRz596lw6Hx7Zudbh1aHa+9bSNtA6dVyAMuHxnYgPKPfUiyb/pQAOpCcrg//B/kzYNPw8t6feh5
TWnodiBNwuXUA7DarB2zJ5h4OkivUa5ox879jj3/IT3UA9eyubTI1AQjBgTxDSsYCgCgQIZCUvlI
UOMp/2vrLTHHC/xiz00YsoTEpCkUX+RX0d+JQ5j+Ivv0nFVSvJpTyb1EuwEOdbmfO3DayZ+oC6Y/
mqmJYxvnzGfo8Y4eSVZ9Q3ncfL5jvEZ7o36yfwjr7f2J54TBTzB/tc5oJV4k4aOFAPc5wsgHUIdF
d6zDfd6a6spsY+NPGXdCiejvANpX9H+BFmWtZ5PE7jhuONEP0A3z1YQ7VyBQpNQuLA8RtxxxoHxx
TEKkK87aSxhlicE8WsBfLznKsFcL/hKXt78HBqRRIIqVh0RpibNVYKD81IvZu6zHMRN4zQxicluQ
ZIFXAQIJ5pIOqikZqA2KWbG/iePPmE3JW5Y4TPEkK0nVb3SOvZgbo9WW2SQFOfbBUrPGDD2O3BZ5
WB5NurF/EhQ6T3nLi4MRZ62Cv5sByK5jyLsW1VVceijHDe0iV7kosq2UIZMZIq1nUMSuTGltm3V9
tOU0oXswbRkfYf9bZ/d4BsvY4PWz3I/oe3XEgchOA8BzO/sguJ9+e/MoTXAhNg2dlOaZ5Ab+fM22
4VBAviCW26H9mrr+QZTsksiCiIkxLoG/DbSkfmr2b2DJbUWSExnANMGxTo3bzLEsvspDFriaC3GJ
YxQtBDdAG+1uSPrEAN3i6LyT92cI8MDNQrV+4DAOAmVwtGT2wQmJHCkc4w+KUstblnKC1ZYOjTDH
F3gwh9D0ZMrF9QqrjCuENOrl9a597t5PGlTq0xzGcXkgGve2TEq2cSx+VCsK1/iYq6jsHepoYvou
kUOTcN8GiVYelP1RQfE440oTXudTmGbMBa8SLpKfXXkj9lKvvf8nvSjb3RDXjhcxZdLPkMDIXv+C
8qs9klhllmiZyzB+fvYubqKJnECyoAdmn5x4fVlvoS3s1xIgXTGEIq35d5/N8IyH46ufBRQlxhJ5
sI+4nJ1brwDV0LkFFFTSeqvU3pi84XihTGRr38ecHyiamTq6b3n7KTXbZfLDB9GoPCVdtLvQ/97c
B9xpc01LdWUPpqktnlSX6HE7MH49tj9ZpJw5MV81+/Fphs2ge8jjZngCDGr6m1mOXmXzZKue80D2
nB/Ez9xfUEZoXpSG0pIv4lIdfeb2Cf4x/NSC3NI+c/5JNS0lcdrm8M2aYRKIaovhS/OmQwMWF86I
LKQQlxzyeI6MeDB1ZX/x9Y8dwkLA+ddbaHYyk3Yrg5KqviDaBoxvyUMXP4IviLPEqXagsyOrYCp/
vEHfMHgZFXcRukCzZvI7hwgpCgBYTOCnpSHK4jWDnqosS29BSpos1I6QJbD0Bov6N85cdT4+I5Hh
oKYphpZs6MS2hQwgJDueMf8ztfICuyoJJ7ZUU7MM09zTrGvHpRJkyGDtV7dsqiWTEgaMYPfvvZ2Z
6jeAWk4o3bn4gcXvg7BsPIwuTSSn5/H2kHi5MuiipMSCkzF7a993GiCu3g0x9JcGRZU5/W6nHdhI
VyA2Rb6GGbLJ33n4MyZt2FKLwJh/Asq9RM2OO+5O0bGK9YhLWOrnU9tsaTFuOtEkF4Vgz/bP8YRT
7YCaoW2CxhEcbSJlov+NTU30blIakl2JbaRmV7PZ9Vgn8fmcsK2aLbLBKfYs/y3WM1qBLWDnP7it
IR7uBOWLsV4r6pKKT+PhenOJZ3s6dH4VEhXZuQ6z1usu2afP09zcrw5DhbGo4jefcixzpnsNSchU
J422Ghouw1HrJmKw+MgLtS1p60D1MHeTkGPqLmbbq4s4vThYmSZFRApVTJbsElNIURV9BX2CxdWr
dYSbQ6viJcEg49goptloOIjwnezF7IPG0eP078q+vTON8oaFizgaXX3dxfNwpcuXXiBMNy/WX9Vq
U7BGWpTVgs0usgkeUbkeY1kVbEPqGYOgPGl2sOGOM6WzeUFBvxjKIxwmY1m0cUeboN0XZE/u37NL
v8zh53XEHqew/kIifaA6Q90yM5XxP9y/JhmzqMfs63IkTHoiEmpXHrgO4T28Ntao+S9aV4cvOUOY
sLPNXef9P+LsggJDMnh3J0GLQMUGR50GTTU+6c2hBusIly+N7kgm4IAYqBvPxClx9bJ4UA9PP6ZA
vOtpfWzoHArtvjGGaddkirQ5EIDhpEb0ALq98BKibWPe2Td5uObwULU4nhKh9rGj3Xq3GRIQcvhn
g2cmVq+fgjte+V1p+nQs+6t4+U1NOdQhg79aIPj3yxit1ra/NDHLgodQ0AQOJ9YPQxNxOvSqSTUC
PGOJVJyF0q4ZI2cCdgv7M/hrtILTtcyLecg6cOd7W3HU3D2mc0hpFe/myguHsC1a8OsN+4g2dQB1
KJ5iZn+ixy/Rm2oL4KC/K94Lxjv0zK73CIHS3r8EL6y36fmBvnc/QpXL9gUJTExUQrle7wUYwEwB
RyYyr99wQTVWPNupPCgCEnYgMRY+rE5fojo7LzJ+GtBV+rS021eoxbknpYlPo3DK7BEqfi3fAGis
FPzgAnzbtQ1ZxoAMjR1Nrg5JBDVvXL4vLVQgSHOQI+OMd5Py2OkB42MdJJJRi8cbCLGKPYO4Hw9w
yaB5hMgzh2wGG+bo3xaJai8gGxm1CapFdBjtgCZJ6xH/Dbkkd99+WIeQIszXdiKypt4HAKSk/3el
IJk3TJyk2hjgQRhW8t+DEU5jHMHz1E/kVZ7GluPTlrGV9l40IjtDqbFlzukBshitoBUYIsJz08Pf
/yDTuLW+vE0UzVhhFOsSWfZ2OLs94OritLtxMYCPxVTHD7YK8/5ZAnEnvmeq0wCmpnna/GeysxrM
81oOhIvYUhqw84FMq9/G92Fmos55rKgXntW/1n57shq0qblidzd8gM0J4LcQWqLpeP9cm8f5EmXO
hn7V0Bk6gHu5wIf+KhDCDaK8BwvFo6hVt327hACaanBQBOJsOgbzMssuHUA8K0tjiHldmfm1Xod7
eMfguOJi/FGg8JYPYWPbxIUQdAvkebTZmuNOq5aW9vLIgKnT6Ypro+/7pa8OFDyV1Yz3Jj/uq8Qx
hC/ymCzeVFWkYwwz5ueweNj3Fk+y+Qof9Eyoph0XQWYPoRVFEe0+NSXxyH/4zG/VLLGBjl1zVv6y
4Iu5BPW0tu3dX1rWHSPahDHexL/yW/d849QII4P82LOcgNniPIR5Mt5a/zyXZx8adYyPjG14d8P9
0O5YJtGHfg4XxGhFjrSMMfERMRSSwU9J/FsnQD96IhUABazPos4Q0KQgGY1gAFWc85iayEAF/PUY
TsYddqNNS8ZxiSZ9wAgPGL74PLZWWGqk9iXBk4nMcAgggy7I/zuGOnW0Ieq7HNf17QMeCiNj81B3
7hCwH++XwGMAsSocoaphN8UciJOojeMDpGcKB/1kBmxJjfKT+e+XRPMbkhHSXBg4553+PK/AjL3k
EbrHMemhw/lo0zE6qvqR3+wYlylyEKTFwtJZ/HGWeMReH6zbd2tXT82AbeqPfeUN297oUORzOnmY
AO1c6jHjmCSxvjB/v2pBQcCWidnM2cZlJsGfDWjKCyVHHa6DHd4yxiRpcexqilcQaAe+fCDwrAJ3
F2BJJAgxhK9p8BRh5BSl44+8bksLaRHyV86XIPyv4R7ZcG8zldGJKZFrOyDWKNhpPbXRIhpJZvVJ
hITYZP9gWSz0BWWBL+4gdVRjognZWsiINCVtoS41pidyNKhu/CTxZjAnwcAVyYythEMBY+wawXn2
CKGnCC0GVcT2MEDkUSji5KwJKcdlBBEcXfpT5G7Xc57/ZalonCYQoMH1Wr1LP5CYbxatnDxIcPyd
FqJuXxOAbhJ0yaPZuNMkohI3m6Xgx05QYO349O39zZWSsvkCuFSFac407mEAYzuD3QpKiriwagGU
mN86PuGrMpZSiVPI3dFsHNeovC37SAcB9yUVb+IS/KCJ2SSMIuGgwiFTYiqZYfENie5h8ijluDqt
7VhXEaO1/zuGYvFjGL9Ij+ZgjL6jRk4/1snyzWpnRn2AN8X6V3/E8BoL3w+C3ScRnAWgu19Nz7P8
dpxbKcc5r3sLPIn5JdW8++LITOaU4fAiATntYoYS89a10wtlbmgeqJ8L0Jv9bqSfaojbzs18LcWM
xsSO0zbWYUMKpPDbBQwV9yN9QeU9xpwF02Jm2sdMM/2zkPqpy+HqJbeoid0safNAZMnOBbQ2q9yk
iVFevPwLVh4afkv+QsBsdNGw31vaHmibiSJguM6RhBv+JsxOYkOeenTK0lBgCZwIZ3BWZ6RgCjRl
RN+BACLGqMsIPPOZ3AsUlqypu2xusWqz3OGHVt2KmP8jYlIE6UtLWCD1xJSggEZl0jWgJ/nWV57e
yIxxQsEqKU7y2Y9x1zhcWvZkX/uXIN5KKrXi69EC8aFIPwsLgP+F/hCyd2aP7DFptq+zVJ/hxgEC
NX0EEa9POAINRpHUWp64liqIe1Tp0oYy06z6FNxJap+gUBKNNLd0dUJlGg05qbHB1xRXTfpBMxxU
i6HuJpFvKejS4hmbztZ9crIh6ABRNo8XwJ2/AHXSQPkC374ZUga3dfU5QEWQrcpUYiFPhJLFJAGe
Y/0RB+T7Lrd4lfa5c6XXZ0eHW3UJFciZ327Eq4hUDCh3JRAyEjPN4OiSwwITpWUjsLlE4QiM+EA3
Vz99FJJCVQjVTpq7PSyjRRCvExF3EkYeJCSvzBJO0gS+8dRW4C9YGi1B+PSZSVpIU4gp8tUEcffy
yh8C6aMc/YgMBPyV8uAZxd3NoR8TWPiK8zrl4Di0/uULuZcjQ7FnQxR6ONLGKTgV4j4jL4Rb+jj2
+4vv7KZ1WNDzvETcoUd6S/+80/aT158K5X5ZbQjXB42vMh+A7ZWksn+Ddiim/jWqiUeVT5q//4Ne
O+QMr/HY7FhKIDA9k+CFalBtV23RwBmLncYpUR9y3yyIuIOcJYWvEqr4+cjOKdK/mxwjape5sjhI
Qm6YK43urM37o/h8XHJ1Y2BxGVkxVoBmQVgJOBcUqqmvgGBlR+JIPLNv+wkTDlRbMylAPGqCDAgs
1ln//+ya35pDV0IhL4v+GWsBHWfvMmTY86Udl7QFIye58qwHOnnLVfpzMR7dZknDiqsuuud2ittv
6DpzYDK92VLeuQm2VmrBv/ACTu6o2dS+V+EyJdU8pupTlgIQIyIZJGeggDljHR3IFzM+Bbcem9Ne
CtZ41vSYPNltKD5EcfgXjiVy0B/xiBfzXmtS1245LQjrZ7WPOgkJ66qvNpcnOuab1bvAm9/jb+kb
UPnfE0EwrvtqYFa3hITUkp9qPOUVY1uxZEW9AebZlxDwEcJp9c36csi41oY+vugQOB4OY6PiVRuq
07EICiETeqv4y7swOSRg8R8rbf2OngCN94+sjojOEbZZkbpb2l9Ix4yJ1dDwKl3DIxyWDObu6sWC
RW6Z6jqYSWXegYR2vXwN8IusKJw+jv7BlWdNwAU6vt5kVPPfpN5RosDAmHB/jS4mYVetcctIisgp
T71pecgN1Nv0Wn5dLeWWoU0PHZth59i+IuyXsEENNy595p7AiKSeNQCHsTUId/PDuKTqWP3bVbPi
Vwku65fHYcZJeawJkswxtmIOpswAiIoVK7ldYTuhv9OeggoEmZGSAGDWpi+uv15VHlJ5ngEXqA0d
jF5Z/AT+DA3DDgAdhN709u+RE0oP32TzB6uXjzMcIeH+D1krlLNq6hO0o8aci8IqB+yW3hHc59OT
qRzoX7k3eyxhqrtIC3c0TMJ8Z0VOq8OrmLMJSg6BYpsdm2xuIQiTRmLCdCvlZMP2AvoJa990BYAN
M+SjFK59JB9jbKCJLDrAhxOyt1HRXP+buA3qgMlmZrjZfTF4UElV37EVnTHbRpIjFgMO/TijGzxR
LrJ8iePEJBZstGzcB8/b/a4VLtq5x/BWy/uih6idrKbgPQfi1bC2oEvZpSOMV5xpRXzMRaYn2Lpp
lg4LV8Nt3KgmFbhCl2ElyNoW/thfziox4YQPj4LsIfCNBTqlIDdHzMOUODvs68rm7G7+6vby2myY
/DY14FyaNeNHgTcHk7dpsRA7YNtcWAPRGprlpWrcu+0W17Cv+uHRWiGa44j5woug/Pk4500hgPkS
01o3XaMAprwp2hEytRlqtJ/2g6+x5jsT9WaMqtQx9JMbOEwMXxdHM4ILq47NhDy20JSyYs/gABBX
X5ijkqGrHznFZxJujAjO98452UZ36unapFiek0Df/n+zxTLivi/xF05UzEzoLqvMpRPRr9SjxSXj
ZR0UFWuG/Pww4b4+V8/3ywIYK3kQjSk4P4BnRuawDKhlTQTK2br6Ekc7naY0T1s60l6iX8cEc0Wc
5TKgOXybASrqMki0xdxF1dNlRD8vo0m5rxLye7KIJ0q9c77Hp15eNkRAGMNfbb66OxokXoq9Kzdc
FF3Hsxhu/n3ZP/iyOY527qYgKEAq30XqWejuGDwhlf3IQ7O+qsFYdj4kQ7ICsh6JHko1pijL5gSO
HTL+N6R4SJ5/GlD+ICE0lHDLNctrga+4Um0wuFXsup9Mzk/qCrIZgWp394Xbw8txx5n3DoE7JAAj
ZHqYhuWAENAFl3tDCUvRkZGjNWB6faIYvicar+xSz+lr50SXkdt6Cao0BQ5insY8KZoxdP6oNY5N
2UJhszk3NwLvikLbHFoY0ZZkNCqZUJKcdrx9H994hZX19j+zcd6ft0Wg6mmPDNA6PZ9r4vi43Z8Z
Ym3JvfXvSRdw9BsPrbIA4RzLouwYK9nxdC0UOL2V1rbFBPQUY4uqaG05WHRNYbYdXqGluJy9vKz9
fEGvLMvKStFcm8T6uDYX93xBUhieDEfijvfRzugwkvFOxAfjb9r5wRm1A35mBjexP0aepIha9Zg1
xdZNn4ceDn0HawMIOAiruwUEoBg177YGOu/mkDyx20iBGXZ1ASHAHcJQX7ZnDKtJA/4EPzFh4SZB
5XHOIF0500+xM6iLoZ3UKI8MKiP3HCq41VOnGs6SK7GCpN10NNLq4fwk9ePbCgxSXpJfX45njFZh
ZzEfk9cIdY+a0G10MeEe5rryW4o/VbI3XrfJ2mGkKMGDh2yORt/iXO8va+dH52kCP+w+lT9oXILA
42JTJU0uaoUwCKWX50PDzyY/dGkr3uAAC804GFlQnRgTAG4/0/LQO2wVGeXpOSSsf2preVkpEqU7
5Jx/WBxvO5ZpITINCA9J6gaE4f12rzu44tUUd3iQjsk/F7iDnqA6y0790cMEJL5/a1Jnmfs/mGIX
X417lKPTx4DvgLm+GepmfWtA9y+NaGgWbgdnf64tG4uq/zG+bM5DK0CJk3gn/BTZoF4yHBZtJOaA
T3SElHfd/GpITx9rfaQzNWwueQoehmHLXd/T846AS9Ba4w2Z5Fk9TRlbuSVb2cy2Z/G6jb7tcAZX
cI0HAtM3xlkKhDH6T4wKlJo9q4+G3py5E3v8wydSlRJbHUrahhq60dmwPCKWcLmQ/T4OKuBMtXRK
cpteZa7yHY7DR2q2AVXoD7I4DaRB/VglubGnGPvcaRtmHi9b80t1I7nT7FqzPHkwW7uhcagyGFKF
2HnX01MU1XlOnwj/EO22Y2O5B5gCC3+ah8Kis1niaalwTbL3vuAuRAd3FgpL+TBgCtYT33PgOQeG
6SdOS8YmGBnlplM9B1PGTAq11TEX4d6mJwYj40AW5eJGMBb1KUX3aZfx0pgk1zverl3T1rBYTdRW
1lrbx6rKgWN54YvvAXAc/CpG7L/zkxKpLS62JYUi/Bb7hlEmGRtv6rnADN6OMUHAlgFDN7zu9+Xe
CKp6YUSa1Te9YyJEX2HgTPxlwtha1u4Hr533461Ve6cXNnpuSBNfedb/YtDZ4kIy4R7zaj1UIssS
cULCF84bt1bnfFTjQkKJpGQCA6Ww6mEqbSf57wv4+h/I+yg9CLO8tUQBR2+AUV103ifYAQPiac7F
kVlI3N/s3XW1S64Ahlpa1VDV37vuk40S99U51wbNJZAe6wlvIKQcK3ulJHG5EAxtP6MXnfODFebW
Hy+E5gVv3g0JaDS3P0Bu/2FPJ9EoePf3R3MIR6Pj6gPNEPZtX1pYe2qOyCMA1BRxWRlAr3X6h6m1
iq4g+2JmOs8sn9AlxMt4R4ewRWYt1qcZMRnh9kCYSkyNCHrdFpt6AObX/PF70GeDgOcpIwel4Z9n
GPP186IqBs2tg5BIsgtHG+LWj2UmS9idV96TQNedx33P7i+NGtYWDQf2OhShQ7/QqPffulbOJ1Fc
eD+3vPbUS2xP/9e1K/5Ayvf/IWQfBnyhHe3Tae9do805HtNwjSduuUd5FLk9FDzWkZK0lWn7Nkpw
PALE3fNfo0w4dCtmZDac1ztFBdumHh1uRXdZeC3cvE2sgb46/pYz7EBcATMOAks8wkrDRauNUJ3H
mb0XjHmTvOXEgrQ8WfyYHwRxjEi3/T5g998v5dA4E20AKKFijX4SXC5EaUlU89SngNKPpsEI7fHu
9oCiFHOzlGmEGsO8zLZp+iB1w5U2T9mFj5nIrCs+zUhgPnFqhdlU4114XrLkjXHigGgMvNBUDlgV
Ulvs4KofIg9bCu4mAP+sX++gDCav0RlvgLH8QGSAxeu7u/Op/ZVbFbHD6K9vfe2UPMLaVOfR6NVF
dkUM1FMnNxSwlDo73jgp0i//0FG3sB8Qm5xKvNcYdluFoYnyrfBgaWu2tpSoi3Sx1981pzXp9sbM
k5i+f8Q/tnSRWYU6/03Yad/sUiCYPTt9BRTupFPmUIJZQcP7/s3HJdu7tbT0kIJ76GSP+2hEvq9s
3H9p3ZCI3FuiW7d/3Lok7oRB+FNJ8LzkK9Kc3a4a0RQCmQQvnPKHJVidOofCvCyxqKHTUjnTKeph
i35g2Xjo6H5/VCumx5WGVHsjdawbp11YR/EE+4R5XEGCr4WUJE/i7td/XvfFBY661Br2vP5aan0S
wmq2g2kAwFPK9h4u4iYPdIoNDe2we6AHgWaTfHvRyCUIFYVWZdnRBwnDCutD/wY+JfPJ5B2nptpJ
LXVg/a7WOSdeBDKQg8D02JYCFTHG4pKFtuCJn71JzxgfB0/QwP6ML4DoxTgGg4rqowsVdWWoBhQ7
5xQdJk7XhTwN2KxiX3kUWrzqhChUskx97qQlftHY/h4Lpeb54eg1SHVHhWwZOq6/Qtk+fBGdV19c
T8OQXVxTNJsBj12/0ifSEMWmqtx0tALgtoj4R4WycXdGFh3xK10fs9yJ0XmRx3gtrjmkvXnyu6zb
hm5B032isbAOvRJBCSoq0s/YRtr05C1SbhG6RfyQJUr8AnwZ+jeky2ZB2nj3xgAhyA/5kqT8+TpI
f/Rra0G85vKjwbKq/1fynqjsBa7fRLx28Py6dgJxLlnxjkEmKFiP/wmzIXiBGU6FCnvnUxYJeRZf
aVCSmV/3NqGr/MGfu9DR9YuD9wUywO/hQGoJfpI++jsneiFnE8bB1st/0fIhdtTlb/RbOvr4bUJg
/myGlYQ3LIU72ZNC4HyDJKTl7bM/vi84hc/iVvRGWi/1TEWerWpu2ULgPY3cBCa324GqlayjArIW
um7wEpeaqwc8CcZGJGuzpFRKWe5qgVwRTqMy+CKueHORH7u11b/hgeMAlMYstHx9HGM9uS4tM3TY
scj+0IwsVsndXOQiMFj2NLpO7eX2kSAjXR4yBCdDK2tOzyaM2LA/erRXUldr+LboDxPBjoEhJsvP
Qf0LzgkCoj+PhdgSJu0hW4sryRxBvxhGNnJh7LsRPkhXelZO6fKZYrfJfZs4I/tB/dtbiMpXcBPh
Nl5J3a6LiXrTCuiqk8vLtG37BXtbnRQF59lWEhO3NxfiGScwesZTi6Mgc2f21tt5l77tzUyosbCP
bw+QrBd/2jnVakHI8VW8OBkTTatUUdTd8DojdPdlcFbAa9FcgR1vCg3fTp5R3P4ukR2z0soi1Xsh
wKkbesjVWuub3s1J5WrPycUn1iuBfTjZThSkxbfVpp4S3F/3Wk48ndWu0/KGbSJ3d6RIWmvhfoY3
7hOphvo12v8ko0s9wHk7guUce7NC5mR313PH/TIh0zmN+pG845SJsOIqgh4NoLDfUIKA8YirUDif
tZpz9u6HxpzfgvNAJ5HLNB3T6s3qPEBDJQ8C9SSv0nqMCc6i0uvIN33S6NURumoi/q5F8G+RXW7i
t3xzdlS39H/9+2XxEQXOoKyk9tUmfP/FRYbvp/K+QeFATWiN/SG7JNcAJdfHg5TZxSNTXjKzRygx
9guq2pVomEVrqFsaoZwPNWxF1nwsxcyHtx06EGw93K6o5rrlr3flSVG5k86NIUZATt4wG9EtghQL
2G2Yw9+Wv5EMD37Nm9ZBKl7pXB+hrRszcc83jFNplWtu1dl7Icr4HHgDe5tPPeXxd5RgzPUOPNGi
epDk4Km6vLnixYuWWhOaN1IgqcfoUxrH+wohsyYKt1gVN0HCkh7rNqHj0UzNS1uA1BeeoENAnUHu
aPro9Xk1MjPxLaP2LLle5DM47fmZ0B0sIykXUoi6COpDUjLNqaNW32f/WSNgaNlZIaVY2ashNKkk
iJKND7p51QtlgRwjVOVUwFDhNX6HO793UgbwW/GaM2loMkHqURobb128E01PoibPNX/zlNtDTNEz
0GCNJR2JO5GhRA4bFeclAM0Q5sXcqJTU2WzjIUZ3vqfA8qS9KXZMF3ro8PTsKi7E5Ur7hQZ9wTFB
qQZRm3fTE0JCaDM+NUC+4YjRzwIOYuhr70M4+CyY3EBjPY5rU30Ef7q72dQLy3jzSuvuutkft99/
jdFhj2nLlUcl3J8tDCNuCrHc3FgrsOiX8TbM2ZEAo3/+ekkS+flNT8wAq0ibkcWycAeIXID8Qen1
tNnTXTCIV8+jsdse0cyESdI9ZBV913YzSg0WwVQIWKVrIPe/jTvrUrxdicF5+1M+/v02Fvh1F6vz
MBFgtoZpw7kRWzZQz5FojMj8fcDZ0RDW7I8n7dU9GQV4aAbHlK2rcTQ12XpaMGpHOm+QBGvPmtGK
houJajOo0DR9RKUJ7cEEn86QbSAHswpdSIK1edw+2dVhyGNeW1wh5iWzFIV177vFe9bMGQAUqsbO
nNNf5tFesJfJIpM3c4Doq0nAQOXp0tMX4dtGXI/02+KkMYc1mJg8zFswBATOSorWVRe1Ca4aoQul
pyAdIrv2P3jJOI674oxPzjg99YhfpZdBSEbmtosHh07h7qW/OZulg/Rf4ZBJzpOcfHVJBZRymx0R
DLGpSTznldXsvrwBIXpPxPn6Sob0hcD+ADV4arEBEkjRi8KOTtuUgY5elu3/4a55ruXjYZ+8hZss
Xme8JVpkbdpjlPWg67t5yrFys+ACN2GunOtU30TMl+T9b6bNXzA6Dwt9nhR/9gVj27vBjZv6fWW5
eciAtkYJYZD5vLEIxlAIUaFr6OcSo0saF9vkxsyzBWqTMAL1H1UiJSPaq5gmr56iMULOvS7GNUQh
nTaWBHmec4G+qRiO6HUBz5EAbuxP0r/+ORkJlpnuieQknoqTpTFzgLkEw7uvt8v17n6VELkZjIpu
ZUd1ZbamOc9p3z2QvC5gVDzjN/BvI1ZfSTN+8ZW602E07wHP10bG+KLyWsK5wQwohBZGHMHPhO4f
K87nSYt1TwzB/Duiza0rU5UxnIvlr6+4RW1KplCzoIoZonbZqJo8OichBhf3OdmuL8wZSszyoF4J
ZK/DcF9jmJmKh0aG1+Xw0PF/6mdJf/hd2Oj5C18zHFNJoey257Pa0+92cpR9bKN51iLYP/qMZ+Tv
Vt1WExl6j7bHGtm1hw0KKXUnh1RiKlFUNBecxwf63hcP8h8Cbn4T4iG4x2TCGxMR5AOJ5g0c6oT3
SDFiWeH2SHVff9oJpa8yVDO8j4VUJz/2OIQKQmZCnwD0jeWS8QnkzmKhCe17q7rWvUKp2DflLlmZ
r3w0+p3Jj8uAGmv69P/Ebb1r5eyLMMaDYapvOk0Bdwm6qmAx4EqBqaGrcxiQEDouS+IGThGOe4b0
K7LVs9inHiRbsNz9C63/a1LK97xswdUCcccSOwvZ41scZq6cd4dvvCjYS1owLDS3pDis4TDIBC5g
DwSkn+py0IbZPK1bO5qCIHP5lhyI5LNHzfeSAuRFCxlUbPmKhpuZ2mIbjLSTsi5INga24qBaOAL8
zwJAgjhb/sUWrBWT/+PorgqDmWu64QXJ1N1wVJk/kiEeM/bKHUvp9tSJnJpTm9JCvGYMVqT2QAN0
qpHxgVHbiX0Yyy0ODM3Dpz31SrhQ5DBb3ktbJhSoSw5tlimn4pG0CFxzqItNBbTfsTsYSWb0iAWk
ZOnDR9OnHXu/mnY5+LHyySYrPBiWPVKV20dFtzpIoLR5h7AvBLOam1uIS2OowLUgGQ2Rr8H9cD94
WVbf85hCtwJE3EcxMBQwUrdcpUXs5vOyTg+DHj2V926yzaynWMpx8F5xvZHZw7L7POi/qoTim9Un
k3R2q4WX3AFaRRO8CikFTO3Lw1ssFo2VOGHpLY4gQZwdnYu0wUf05vkS53DQJacJZ6VOP/Ly3L+A
dzPt+PXXvYP+E9mh4vwLJuv4vtA6F5stoReFi7gtcxTw1nbuV8gcTW0/5AOrY3nB6ZtqIDg1LJ1d
oVeowyilKoLvBC/rLh/5Uaf0Yz0Wkp7NOROuyCeSdfvudpaa+eTBOfRA5HeH4a/uqsqBkvvHUlPH
lEp4RgdgFd4jH2ztQit8P4fRcjf/xOYd3NRav51C4cF+53YisOuWBCUcdPkzbsixa+Bkrd5isn/h
uYxch/lHGBIFDIsxvrGdtbTRU2C0DCZwJNKq1K9wvoSzfiJ1wPVT664OsfJBvyi4Rz0N2jYxpXau
eHvOAis+8a30SC49OH9/9W8msbBRbU6vzfSNLKPncbufTV+BRurm7Y4U3XJKiWlZPK8oUi7KU7C9
y7N8I13/V0xC5tGymK3LBXey5nXJvK+9X99scAKCnxxk59/R+yp7crFOq+EsfqwC9JvhPkCap61j
PfUFAFT8icPQR9HQyqZMxlDrlH1nZJKT5OWxrt8u9YNMs+etTq0IW2+2LCcKK3YipTu2hvQx6Pgz
daVscKvHaU2BZzIc9+nMAqafv5kPyDr+l/rHLJ58C6cO/dyf9iX8VhmlhePdPmGGphsLhEEpCra3
urCijQTVX2kR8oNt5q2DYqe7PD9alEFiAN0sKQW/WHl8bn4vC1a17ffRtxwXVWwQ0BnV/WNeM9DE
PA/TU/b+jeZrjTVSjj1c5Fso4DQlZtHEZVzx2l9GPsBWEdfnCaWzLKPX4TOsq6tyOPlK/X+XoBEG
DiKYqk9CW7IvTGJf9WWACPc56OLYP/kZ6r+N9jW/Z+yqwfr3zxLMHL/nJs4AlGtv1j1z50yJxz3q
yoVhj5vdcmYLzDE0LvAJdGN+ZP89Ng+wYSNEgax6DyO+wgbzwMo4EoI1e2GpbdqMe9/JXpKVVmj/
H7fVsZw/RvFH2qdkl6QDBvo18cJzc7qSBv6+pS8ikEpafutKNbiAUMRHasp2ln7UjoMv81xnZnUp
U9YYDwj4XWx0pqgid6il3s67A8KUNehJ7B1tiLsWE8rMQocA0WVrzib/Z09Q0YB52Lgyaj29KYaJ
EhL+444KOyD1R9sQbhJ8G1KuWoUrj0iwrf164Np4b9nmeKGPr1ms5uwiJB6W236a3g5tMT9IT0DU
4pRhefFmlEJQkflx+jAfCeJu0kTxf86nfsBX5/F4fXXeqYRABk7d/mjz4cfVZ17mohxW5gNmXihA
UltKuduLzJXqwoqonaHW7vyaLxEAS7MrtO4SqYnxcJ1DnGrmgMvj2FhUNdghWFNlFOJ30u5CpxmC
Fx2fp7thlpGUENbDoZuEPsrGs1evNg4ixjmxokmdfIxT//ZFR3kH3pZBTmafDqXjFgWayqxM03ge
EG2Lg0M7FRR6MwG5Y10c3rrXita+Zk60KvjDJ7MVwIpJXNlL7gdAdEh4nC29bUOrABzhnX4ETveg
s1hTiJ8d+7I/Oo/HzP7k81g1tpmklPfH6ndO/covCQgMAqn/TGICtkpwRX1p9YCIRMqrBfWleh+Z
LuoRpyOEnRxufv4IkJdFbuKDOjVGHS0MNiHFTIgv7R+JMtIFJ8WWmbxQy+D7+DYXhgw8Mnd8Zleu
oFIiqdO96DQCOexKPeJYYXeLkatyBr0QmllE18N3rCJNHNZsdA5PLCERANURzs1FAL13tzAXzUjA
CwVwxnfaTZaM8OFWA+qesMtZC9+w0FS5BI7GzqQdN1aZjZJSTa0y4W+oG260l8S3+5ZMWVOkHzjL
DptLowNFJZifUHoKOzFpUqWy7XPYOL3nFO4XXm+PURYw49hl3A3cCDGv+4ki/GyX0waLRm7sd7LV
r8QWQC+2kqc0qZwv5Sxm55+yj8GUbCiFy1X8h4XtA55/vDKb3Y5uzk/zPebnHt2Wd+OsGFmW9GEV
y2xFFAOzEfTaPuO1NuVuVb8AxL+doawUT9dkG5THO3WMFo5yqk2MIsM1xpLZ7KHCQ4vdlT5uQtfa
2T1JdcKnYrhx2Nrqqemfj6OvxQtLtuxdou1Kvgp/nxhyYFQ5hDu5J5sgEfXlx3hXOB+UZ5OjWAN8
GazG7AUEVxAymwafHx8WbftZ4SAX9RjAgfyHQAo/rDXkQrkEuj7vJgsYG7AUayw3nJmaknBZPf9/
lYjcPzkdg2TmLoHoVuj9pCNOgOT3Idu2+0QBgyduW0Hfezj5rhrTKLEvzddJ2e/ejNru9YyMKlR0
HLJg1sgRWRPTnTRcb6OIbuCec8QzAEVGKABbVoe4chozqnFbiFFQW0cLL5adCSPi2gp3o/Pv/MQx
3iG+uYyuJ+Y2zn6OqxDEKpF99Ci37QU2ZXbgm3H+5P7rxpeJg8tpyobaOK0muuCiG8FxH08hWcYw
aUTD+4Z0VRm/0tTRiDXxcnvkx2nVLZzZOq5XuJ2eTW8+kJZaDGuNwmvJmMrCR14LcXSqzBjHzu9x
Oe6W3xkmid+YkvHgF7wquwOPaZBUWcvgarEGfxG7AZ79qrdxmDPYneb2cjA+07vbZnqGpeBz9eFl
uKHlu83l2XCNYdjVigpK01t2UOPeoKieuKGSZf/JSSCqms63YuRAfH+iHuBbJdfjiqxpiGy+Qs9G
MLjF1p7iN2DG2GHyjQFtvZDKHVRqAOdsl8NoLPzUSCph4CnFtpdatoMAAjwQITHj4J+ZA7uPcHgX
YAxb214LmUOYRuj5ONx5cCuSeUdtNw+/2i8UJSJ8D1tBzmLaz9H58O4qfzxhXoVNq/WeXNF3Y4wf
iZvHBEWcJ7s6FIene/hcNlI18eDmt+dxZCJo2niOrFTtrTnBDhfDr5cRHseXTVn//wdag2P4gGJN
8V99uPVQ1QsauoI6Ayllkf6D98iJQFRBgoR3i+o9OyHYvMM8bv5STa1oTXboFgM2dO1+zemRPaZI
ZZL/vqmpZdKyvPQTlW3meLT6FwVP0VypYTIFlxAFDsoc+zGNNOuxE3TBfUJqvx+VLIHiKV6Nf93x
imme/jB/vUXQe7zY69F5tXxaxxAVl9ZspFFcFUHHC17id84KlHdxL3M+DhOJmoiCAagyP2ql6pEw
kNbZ15GDNs9rj9KzDOEoGZ90cW+0Z3RK7XsZSDWwNxKGtiq8b+rRF4lFWIDpRibuPxAvpCDPAv8Y
vsyYLtAVwd+Vba475QWLf4RvHNnoCJE0EAx99h70OZP5ORGrTp5Um4qq3YCKuV0McP/bia8nOv5S
ZEcX8E1jxF1WJyXSmX2VDWwOD1JYZq+aY8cRvCat4FDCvtjzuj1u78LnGajMXKe4fN+/KECZbue1
mpDAFeXqQeArERA9bwc9ive/t7fHG9QhOu4rhsznRwHgQgNg/G/814FC1V0P1pE0oNbIkHMuZSHI
lsZGtjoKYF/Q7pqnXLWWDLGFLgIs2kA94hwv/e37y5o0wsRlDqZWY8AMCdVAB4+MY1Vg64XLqt2G
YG3x6jWwRzTbpM21j1+Vg7zG4WsAoMfMzHq5SsStza56ixKymLM88r4rJM+/LBX4/5F8htjevHhP
DNqGia4u9VXiWzffcCM7PmZIegp2atrz1RzLRQq+U+qO8QD5PD2BMx78GtvzBl3oQG1HWC+LjZTW
S2pC2dc1RcP8Wzq36Mgr77WDwNpRVG+OIgamrDnWMxpK5ECZu6S15afTsR2qBJ0RZ2O0ycK+eYBR
sjKXTAK6nH72DFoIbkz+sV2isSb6na27f3yQdzDI2SzHPuwCnTH4tK6Lv/+izyatgrjTYhGCBfhF
MkvEVBq0h1WWuOXdY0cQr6UytXWSB2S0TRd2nOMwruYXXD64UDZ0tASxz/OYFj7Hd/NixdGps273
xzs4qtXyh3An7ORoV21gDx5rMxqUC9X7DU1ogWF0SfcnCQseZTjjBjoOFcBgGiL4G++wYya4FHem
XSX+OwmO9V1v/oLufb9zZylbT4ey99RgpltrUkUwos4X0oED/zDDvYSyLmOhvfdWcLZX8KbukQyQ
6JREvvmV4T5g2FoCVs00hDGDbxNsTnil8Fuy+OL2JlwkafzdbBoJJ+a8pjyOZ7iUvaoqkFlSw2ZX
qQOZLWOKt57II0AD8tqugrMhN5JgBS9N3QPFsASGsJce0EG8f+XjAo3rPCVPMZfqcYm5xaq2mJVh
MseDZG6/qn+IIAv2JYj35DvViU6RoQR3crgBQJEZNrp6xe8WncKuR/EZtvtMfcPB/tFWqhJTwCpM
7wqRXwVEJH8BWgtWaSDUP5IHlgIBwkMQNDe8DmKmWhuyl48iYi0RUJHoV2ObgU1PfIT8bZYIDPiD
ACRNHWG2oUT0rbUv4h5WtuM6ToYAc5ITEvEehkL7kg7mbgIQHKMqfvY4uKo7SofwtHAMAN7UotM0
vyGp0YbbPX5U5KzQGdHAnKvIkkUmMmLPg7ccGAdjgGsUo5DaVlwtsoOYdoT1l40OY4OjakxpQ+49
jvT/CeyQYT56bHS3KuZktAVMNdZ4JHN9Av0rLtcj0ytR2qqVLpA76kUIN3kwXhMEGf99cMBKYr36
DMayeGRV/EHlSxE6MEEkmBNDL2oTitwpij0hWghEB7ITEu2yZLOd5AgcWXtA9K+x9k+LnQyyCNiq
N0BklkK+Jh5BHXIwf2McnB0AnD2VebFAJOchzr5uuGbpfD/JAgbM8aYzNOazRW2g/uaf+JpTl0jD
x/yt8Ixwgr0Mundy6r+P39OsEQhCn6FdPorHikUpr4Bp9Cal2VDmh4xkgkDQqTFToKWDTMZIDMTA
XsekjsPJ31dN1QM92IcWGNeJsZi/5CN/SEsZQnQP70x1NORiPPjy995Wq7p8aPc8fNbWiGPjG7rN
ZIr4SjrCufDr5U+qMHI+KeoJex/w1n7zNpKyDGBb0nhXge8mRkPRGYO1uRC/IqdWMCkLB7xPdTly
I7erQbxfR0zKUJGyRyZARZavc17d+qGRN2Rlmc6I+5k9eXWtw+kTxzWeEN1ZOsK0sOtTBZ+rp+Up
vcAeyO4EU/JURXXWyfJEn3QiirKxY16ctTK34FV+/VYGjxXQBQJVawF8eLnbnPqp93AseCqcisBK
b4GLxH854OjKoZ9KlmhWErLKpFSofg/z3mbxIZFj8c0bPnw51Cmh7eAq10y8Dleod4PR6I3KjlLH
Yx6m9Hynf8RsK/gAYdHDOTm/0v7r7P7fQTlURmhP54em0rB8ISa28ZabZHnOmsw3eRAw/1fIbenp
iVkAHlsY05Dgj08MvB7zBMcLNCUk+gh5UHeGRB+YczHJd50dNRTgua7vXGAGInTKLFja+RMFTX2p
fsjo25A2wvH4VVE+fQQ378KbT0LReBjZ0zBSKQin5JizboB1fJZ1b0n+uih9q33e50FFPxFPqO0M
S8xX9TKwjOqp1BacisYSkO/NSQ2vA8Tzhl3uuuPJT4hsGDAVlrbLtCyoE1mVinbrOdb1l/0dWdKb
BBLcGjUXl6F87n2Tez0DloSxpVlc69rLffc1zGsbnYrGza3t941rCbngabR9QeFdX31gJQaRAO+V
zjfm7yiYu91DnpL+7/nAJ42J9m1tzm/zi972zBQWImhwn9ruAh0Kt32t22Ad/o63If1wvjsUvPcY
CTrt5ujiD5J0cYdt9R/FBEO9HomjY/oxqpqCCsyW0Ag93BfSwfy1J7wlnvYXSchqWNcovOrPI1m2
+Hn9sb0Wt53izB3wZyXGI1x/LPi2QbpNHkbeygU8fDkwo07GUCdbOM45on5A9h4p4ivsjmGgjqfb
dJNGyVMk2Rvq8n9tI+qBwqoroJ0Cn+niG2hlcrhlrPTP51SMnvFdYlCr5/aYhXjxOsA/sKF/HSLg
bIkXHlrKEHLRNVWFyT8YUt35b9mhRz7R7dOTsV9O94piYzkyDf+mP516AAy8NxQ01eVstLJYkkGK
ZpqFObTr7f3cipH4y78bqTEM4+cxRSm7LQjNWKOss6Xvs5AvJpfMs7dSbZDnRNQLswdjDyYpoMZh
W5My5KvuUJcYxQY+XDSr6yaJdIQ0u4YdzhXTw3R2lRV/yfP7brpFfkXJtbUmBTB1rj/lIxeR4/RV
yRUB6mtays/ZX2aEvcNKHS8ZFEqwv/3NsT4hhuwQ9m2FfFJYlW3FIyLCPjHgOLVvHNhgQKcdxgHA
xQVBhNAV8teqe7p5AnlF+xG8lKJYKo7Gte/yM7YUK/NNqDEeWe7ThUDjUTJSBIlCADzL/XkJSkIC
ub4LDDEr68AneVstztyqoHENgkV1aT2UMSRxQznXzVo/fyMbH9JTu/7kE4GUwPeDawfDQup/tU6b
JfSbIzSR18LfGb9fQVC/y0Jxt1OXO4ponY3AyB8LlrJAMV4k4LnzM16sxwdrrFa8AAZNfcwq8rCU
7GPqNXUKGhmpO6QgwDZ3KWtKhif1GZoSHs6ScrYedekYUEllYhYdu0/ACXAtgOTuI1RJpY04LRny
jYhheDBh0+LDejHxz89oNk9zp8UIYZuYMGO3wnkqKG8kAuOi+ai+2gRObNDR3AuvKJAUS1cKG3sR
2fNj75NnEcwAPhEB+4llm8DP8uxe3zyX20ev1htlB5DDOiMYUE9/QAIgmQSij8YhoW5wnrMC8jV8
jZNgDgCnJU8g8OKwFzVYzflwtogH+wt8vsetepbFy7DDhvlXgEPbhPaIVR8AgDNIHslUHOR22oPo
zII7FL5C6NJ8sRH4vKhGJZpB/lUuuOpP9rvN7sPCT/G8h2aogW/udpg7XHa/zr+BY9Bd0aOSxfED
wESmTM3pVKa7AzuBCHyvpW3zPNM8ug7PTxBNrfFNAVHE7uR0x8SOPBvdrFR+ImoV0D9oLLgATl2V
KUA4XRiuGiR1oGfLLAAXqAShdozWr0me/m3RzGTsbTAsfYBD3qSsx9VKjcPjTk4Fuce4UwvSTfZF
t/ULI0+NGZPoST0wybeCB3kDL82Wk6y66r6NaNUv5qMv2nEGKRYwW8T/r1lggEpVKhgo4/aIjMjR
UrIhCKevXS4fg/D/wd7CTvE78XwTuNJu+37NvcAneXUJJKyv+sCRL0l8Y3v9KiNClfsCxJVmnn0o
HSXpRZX/hGDLFt29fcal/Uwwnve2tGPbcParJZvvHCBzG87DRY6ELiTgoApxI1QNSb43jQ/P2lb5
eSd1pjxI04x1sBrPgDYOMSDUnToXTST5joZIjKxFcXSC0wgZ5ES8EeJT1Bnq31isz7Nijz1tM6P5
27huJDIYKV28girZJ+L/w2pkv/s1ztT9oYtpC/PNVnwKcJKRcTvoNmp8H+ae1WyxNmwZpoak/0zY
+fEIKmcJHGgePBCureIIshrRJBkw1Lx2FLITUmc/DBOMNWC6W8iP7gCH4+F3xXK14dxFFvzV36Rj
iMqpMcGd8/UgrpCPja0ePXYtF8h2POnZ1dD4QTGUPXeJSWoo7j+qo97KUg+7x9/cP/yD+QS78IvF
OD6aLDP1nNhg+vEggmnylM149C5d2GaQtA/YIoXZA5J9TjL933CsP2bcAO1+jJjj409SWPAAExZh
O4uMIJBFtAsjMBLF36BxNqA+OFtGc08N2daFpUn7orZF/ykT9J9KpBvH6w1+6DZOaZnxH7+R7yEy
HfmkB8T6eb08krFPzQGTTjLmqKrts03wQblkWD2VZMsY7ieGLoVgWNDcf4dhpq8O002dC1mhGADV
bKRQ4oucuoZpjLoltS2S1vJ8qDjiBBpwfd8pBdGRjEMSYJhQ3Dpe0KiHpywD+ivy6bH2Qk6OSvL4
y7BiyiMZj6CPXE8HrnKAcAaBlRNRnq7aD2QjOk1DVF/NwSgn80laJARb0R6Wt4gsMFBlwQv837TQ
G+sW9xOmxDxhItiwepvrtf+W3At0euNrs/H2hqB+m1LUHrbt8n3IO5Pbf7ufFIKrXsaJOrNg6/hX
eUodAUKIcZR7ioUWsDgLeR6vLUm8LFw79FOWH4fz6Cw5GefTIu+RMO5gpgoMOhWWmSTpXw2nXYwm
tWz/hX5gXc/zdX1hIKvev0l5uQmFeWGqO5CPtYJ8PxlFl6yeAG+6JcjdCZryKZWcetZxmq71/EcN
OV2Rlek81R3Q9TN9cHMsN7rZuWIuiKLapzvsjDajFSmPRaJ5GODWjVnD8YDdvjfgLWNHOeBBQJkB
MgcyacK3RlgkZmV+mxo0quGXu8WlERw2+/xPhyiUTnxF1oQ5tHoQY71dhGH87lRa83eWv9+oVZmK
bcs9ru7dM6ESaH2IOoblYyCOkQXkA9H3jKyaHGCUO5osDWXsU1pnISNqCJVzjguq8y6hxuZvvphv
wOIsC/D6Zp3w90ZaeCWIBwCSjcR42bIQWxLhEf0Xl8lNIDQ1rAHGik6JE55LCt1OgC6p0AknzYjm
k4Ks+fQzlmcF6I6IyThf0ISOgkFOAqaUw0b0Mny8swCvRdRbG5wes0IhDD+Bj2upA05oNxPy9eNe
p9HtF7fjVYWyBqxH1XJJc8Kb+8If3ymo26MCZtFXvPNUs6h+QrpR0Imgt8wGTt4OhAVN8VnYA8mq
rnDu6WalZ8clp3/4z1I9/g4FONFal9L6Jk2vGX6g64U/qObHsllG95iuMS1Okzg3sJxPOKFwdIXs
dvt4pn7Al5YH961mY1zPpM4ljjEH+0n1pVnuTeESN0fcKgwGAERx9Ci773pu4o3Uqu0ltNlkFltt
qA+sU2R3O2cktgqfqWxPW6M12Wq1Voqt+0HpTiSGoahcTEBT97oUJmMIzMD5o0dT35FRCa8VvtC9
AwjG6CmeBTdSzGShB3A0ROs0IAAdrQgk7SyeBxT5aXG75UvhCu3YlmDyKsfkFAqJve8fNqVVZMEE
aHnBn2Lrl5w1tGAa60TiRZSvDAsT3+d9KJdRiH7dfttu6J6NP0LQbu9bIIs/5HMF/6Eno/Nv+V+L
4D5ZE5lmOqO/gywuSCUn66n8fqyx8pozOL+NIgCKrwDbCPlK16QjfCmV5ZLC35SzO1/0PB6fIQYq
E+mKXWseDiMGQi2d/6b27V8rFOiXtwFu8vZ8onftlPnh/ImwIkDgzwH+6hJ216kAgomXxkuMLDxB
hzYO7iEOVinX8ndU6stnGdN+D5GaWJNK/ekBrK+z6H2MA4Dy6U+nMDgSHszgzLEVgMzfJ4/sQfQG
uqZvhG1PqoYY2SmCYnp4+0NG8+YoSFTEifcxv2O4Lx3tdlaBq4g/ivxXiqZ2mUa31U9GPhOtDtCB
QNSLhrS/eLenIl4Wp2IfQg6GphJFM44gtdtZyxtQtefp6KDsVMnIcLASETZDor3agGXJMGlFhKbq
P4sEnAbgOJEGaxW5ernOKff16Lgamr6WKGdmmXEboSxH1jlZlprB9yJPeaK3x6dXsK5ouRkW9u0l
jnBDTgvF4TKjK624SM+kR77d7o+5Nk81gHSDww3n4tokpP7S+j1m5gkLYInIpsoI3p9TeCqtS0R/
6SotT4w7eu3pP7vPy+o4WUDxQ4zbKqzhZYp9+FmsgsndJwQzyENFFni0fXQ1Jf4VSt1IhL48nGow
IhvbCZg7NP+Lsf+Ne/BDh7Z/gP8wXPFktvE2Scm6l06lU22bdOmsMpaJVSNyCaqk/4cqav6Hd0Zf
TAMOQso7X3ZNoFRRABTvqoEzi7eouigKZ72rYulhuU/qOXnASxO0PVaNQvZTZ2rcRDKB64U11xMQ
gkyFpsV94tB04UaltQQt1x0iLB2e6GNZU98O7hTORVOn5F4ZvtUy0wHtZj9DhmQy5p1TL3p94rFT
YC9EJ0fdgUm05EqdLD2o5JT/hKTwTIz3EFGzqdjzJrnW7tqOKeSNvkm3uG7N6FOtV1+Eb23iXcck
8o/or1XqaDqzuoR3omc3OMMxZPzH5zwu361tn0PqcdzC1xZh449c1LDVRuE8qLRDkrg2vY/CKBiO
rhRjjJutzvKbb5+XYnvOjkeOvMi2afgIPohx5cxYbNBgmRKQMAe4fE1GWTTR55tPNpYT9bCXUEcD
eU/l/523+8QO4L9KJe7yjj/EhxXzO68AEmNwT/sCbkNS0cMx3W9ADNMd7LRc8cfYA1ABa+MezYlU
Ll+sb0MZRpsQ0rqONaqg2D0N+4rD9QKVn61g8VBQUhHgbjrNJJVIrkbMDDaNU2EMGTq98CXRQtVL
WFhIY6lodPPWq9CKJu1Qb5P70i+md0HKazrX8dG1OtmHblZ95m03pDGu6rblFhFxAImc4p8uFkNB
ZFWMg/eAHniBmv0HnrLZiOztqvQIxIQuY+Y9FU6CUW4rcSxVMABwKNwUoHwRS2If834WPsXfdnLm
wajQYMuTUXpGnNWKbPm8Hu8WyIsOLZkBYFubgneMRhwotK7EtxwuveFEm4l950g/Ewdodmb2NWC6
HNnUf4XhFKqqUWfQlR/jFiel1KBKGkPDY6EFUO93fOi9lN7hd2qghV/ESFHLPyjakPVV5dgPPiev
xlAKXE+ZFQjUJhtcfkwwOGH95XDTOD+TqlvXI09slx+vHYZ9by1J29+EtUXqjvMitzU1QHK6Fanc
nD7xJpevR5CzpvgbajiynAQ0tjDwirr1vJqb5jcn+Rj+dOIlXu+XuUxvteH7H8sXPyDkPSAKLn2b
haeo4qAVScJalhRjiQYG/jQeXtFqT1wqSO/p1D9q/FNaiw5R0ztPvlrbQMKeRMkTbYEuA2VVMQXZ
ZFsWn7APKsr0lZMsDZz/GNXuX+QM8NGQ55zyEwcxjtJ/dyl5zOog4u1+JZLwpL5MiLF98mQ0Ccbc
3pHEAYgPhswPAwryFI7exfeCicI7yCEubNBGORIO2rjpkQRb/3KORjiCwUVBYsGskDGGDJCX6+Ws
DaaXQH8Ffw65aV3m09HuXf0PQMPjxROl+6uGad8Qte9xvsejinDg/McjFSbdvHI7HeACzkOYKxJr
lbcQqR+Y8i9b+UbJcAxUYG10Bca9ZpK4MqZrpVJs9M/uGy/tYuLbTwdCxr7TMIRaimBGOjgyt4cE
2huPTV9R1xoYk4Rzzn94S5x7/H36lBD4z2b1V2pk75PMT39izKBbYD1xwl7Fe6lHjpeQR5NUSo0o
NaDH4GkqookEFq6v4UBVCRxK2a+951/DvtVdFQE8YkNP4wMI0eJw+1f3ibDqp1UgNecl76aKCf6r
0qVGG0Ataswjnbr2/9MdB5Z31WG6U74i+zLIo0dVfhQISQLt7IkGgiVd6cvGT1RF7+v6W2TX05fm
esdxBKkk8+e5Dk7GicrK/2Hjjde67g5SKYskXofdjW7eqKHF2MZ6CBlaVMVQ+vf74eVIlpNuv6Pb
7WC5KrQLBVWKINKYVRTwC591KNUxRILU00XXxf+SCK/z5TeuZxLZP/8Blp8147uDXJAQXP/x4f4y
TpsGYoS2OLaSgy8nKAQehIV9ePGnmbMkbeknWq66sAC2H3+QDflNvrsZx1ccXmU/FF+lDE3SGeeO
DtEdQBTFC80l+Wmm2SmLbLiOlRp8fhQRNA3+sNdZl5TIFSAKwo0rqP3mrZI/mIuSxeqMupEa59Pl
cTWx+Heic/NywOVXl8EIRjoE1EB2wdSuM+ykXpUVHWqod2ic9L5RlJYGjaBmjhAwZx3kbAyEjjze
isGXtvxO9pJR+ASxvL0EE9+wpKA2q7nsmIIJiQHalkNv9OMPnOu6bfUB2SRgGwDci3Ix70/cOmbV
JGdo5KsBGy1vKUQGtY9vb4v848iYRIBANR+kIxdqeSXsbEUo/fESw8w+tdYJMC+rqhZbA33Wp09L
mfKc4/naTPg/XR9g5AcMqCQyQ/K58eSbtKaSa0PWWH58lit2InGAb3rowsgh/wOenzlsA0rS2Qxh
APsYfCyNBpVHzpMDlgIkJwJaQ6oLZnhwTERK+wOYNR30Q332miR+Ex1lOi79Tn9SXV38TqEfn+zy
+FKjCFGsBz/JhzXd6taLvvHiThosueMHJxvCWtDD6yXMFRCjkbRaU/nufcplURIfLMEUkgOZOgE7
nADZHLPV9SdBdoxgrxpyKAmccEqD/ocshBZFlr6YXQFaigTtRSwQ60bPhyIJRDDsNSad1sZ24gVV
KASHgh7KqwdaLKryIzdGbRsuaqPKPhI7DxK0CNvRduVHkJor3tkiRPTe2kkTFZ5nmjQot5uVQQca
iA+MMcHbmcJnUG8b0RzNEG6THteMW4M2EljZV3qSLz1Zdhpy1HWcAo2SqKgnKkxXO4+4Uhcst7aI
wYpmazgzLVACI+LBwjD91SD3zAIi3mNsjXz/+pjtpjk1V0SGdjrvh+MFVoFlCcohGuI4tW9P3KdY
qtjlR63cwf6GruQCz0JNhVCXJQVRaq+XTeeLZUMjh1GLRhjBH0sgOQxi2/VnUjwcc4H0H+XqCp6+
CkyB4Mz21CtRhDXclfocF+nPlKxUHysh44FVb/dd3LAPbA5vcHJGdVI+SMs8tYhZDkRtSqRALQqf
wToLTTw+n2dAgUspD8Atmq2LuSQ7GKYFJC1DRQcJ4U9WGLPrxROybLG0ypd9dZ1znOGATAfNx40D
zJ74te8YvpoyNVwaMYrS2GeFD822rNfaaL/ISe4YxbaHNvancqefV2cMq35qmQChaQO8qfuiXkJ7
kWczwinPn+FlVzazd3CcgeaBfa2/ySkIaJzGcpB1ekuXlt4g8ct4niHcyEXLOltdotdmM2Nbk7Lv
YfWHOR2pIQJ/RYTEqPj60rQJHX3wkFUWlIUbt+m/BoslfyG/vlxBA/wlSIIxKNG2SOY+A/X7/i+a
xbDqACMIDOS/glu2tbQtSFSYuvFmSMg1bC+ZmUt3BlHFNHKRDZOAUPvbQ4tSQFYKFiOkTO/fekdG
0RS8FUTlBJlWh4HZ5gDzbO+fnSrigjazdiAnxDChJRAPuZSxFqXPqK7MiI4onChQDJqSNPi+7V5M
b9URLeGGgg==
`protect end_protected
