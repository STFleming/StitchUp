`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hGfDac+z4rHZPk9EYeUjoovVNlwBAyAj7Yh6TngoghCfSl/z+lEiz7O0OBVlByZpPFR01+YWyEoo
QDkBpej9jA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CM0KuuduvZbiZ4JXrLcuhhXPA3x6HyOcpomZel8HI5UO9XFoNvWJtSFltmrTvr2rWN3Fz0qQsLE4
WfUSZoRygtwy+6zZ6DpWOQdY+GuzXffBUkPZCgtuZdFOuQlLD9iX11p9BO5hh30AcVp7V2h+1a5l
2H+n58EQdPqqKI1XiLQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sLPwGO5NqFf+F6cEF2V0/9de/Psridm8Yp91tJXXpYBav+TnZcKp3f1oVwCHfSqxESoNtUDw3BIw
NCyaXu2Qt1IdeiuczsqSPWrWZXmJ1kyJy/CTq32MdTDlsok5iIkqo/1mMocASVFJjPL1INccHeZ0
0z6+hGXlvV3BK9JO9qtlqE2PFu9dH6/IF42J0Ewim+Uygx7u4x17JpK37AkUpPGvX3bJQOE9kiWT
6Vdi4c2AaLTqVQucg/jD2ol+QHUlfxxcjlW4CVLAypMiBTfJ8k8DjLc0rmMIoR3Bh+11q1Wj1F8W
ydgjKr+/sCDngaiu6PbvhmG/sec72HzoGPY5xw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UMO3iDRQXy4EYiJwyD6E1/VVwrmPyXeyFn3sHNJSPGY5d0O3dd/bR/g/H+qhuektH/CsUqxFrPsI
KupPFPmLN872AELCTQ1BPnFp7aba2v5QTo1IjrNU8F1U/ekPwQbM1RtSaHhqZqDLozVLQgEL4NKW
l+TYGdTmBzfjMQVW3TY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Pfh4qTD/ydyNlT4iZ8adWbgQNwefoxv8h5j57xyDgM8MXm06sxxq8hJcJhkgPso3YnUmyN18zc4y
oEpfMyZqkgMzlNgzkZ36H+RoKTozRhrKN2X/Isgm9vrev5c9luwUhLKrda6BsNtwIT0ri7/6/jFA
WiB/3FPAZ/OYsimQwZuTzMFmP026uWW0/ifkbsY6EBbgK25WUMVdONOUcCLuzkgw4HVKiz+PRbRX
Qjlm1tHNM5vyTIBC2ji8MV5KR1tasS700Ff4eloYX/v2+XCXVbm1TyjjZEzBDfF3K1HjW8GHEBK0
VRZ9hu9nGZShwAD8y2x1RgeSpFDlRbHu0BJ56g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10752)
`protect data_block
T2a7picBhtTZ+l/KjhB++iCDJ2DYJp5E5zO/4yRYqV0pGAdCO4S/1JcUQ/8PQMaTUrCRU+DUBa8j
wI2akKMIed/fEDNogDpgiWxlQRX0LQD4rrdcqAxp/CmvWk0gTzGWEMUOkduhouxBslSPI+G4KP61
jQ5T7rLpv9i5N0XEOABTk/CZlbhmWIS0PpIABSQuhVVPbZ8a98y89y9+oH8UGfbEqIkxj35IY8Is
fBioe/yYO8LAHc+DZ4KU7tbsaX00W4YT5qHNptWtGRINCNNQaQWzZ3eWfYqnf3jUU2JHDBw+MoUt
dxO+3tgm+W9j46QQgAPqHwoghDFQM1/3/MJSIEIC6zhQZwC1vIX4eG2MQDgi+NnpU1FdEd5tctKU
DMcC3XzRFSFQfiOkvRVeorLcyrY3hOEmXRNyoeFYvbaOA1E/1aJlomVMrj580Znpjfjbn6xowAj3
qkGMm0p7KFwW27gOsbTNKDN292l0R29VehzAnXTT6K1IxLMjYIP7Pu8nQGdhG7IFSHzfecge39Sb
WXxNKvZd9j/2Hg4yDJHHxfNrcJHu2aBYLadsvZkbDlHMLMJ6zZt5m8eoIFHT1j+IGWPwOZi80Sij
RckQRzilfiZRn6SIsVRleEtjHZPELlyVcb6UdBhHDfdBkWgmK0JUCxuXR/28JueSv/WPdbbA2ffV
BQSDuFSDDLicBrVRAlY23+GExoo+n61qhPlMSFP3fsU2hmXDTQKJXlwHHXl7501RDDw69h4RI7zq
hz99Y+P5AqJzAVHQ4PWmERskAAA+iM6IGozxktGxkhcpFScCOFl5TnTh+j8mudw3IGFWRAq0ARPd
ccVzWLxjHsjdVDQsEgQcOdoBOF1b3wSf3PjUzW3YogM1DkIvvXTvMCXXyJKiR8c7vUyUMacz6z+2
kPS2NpMEo3paGR2Kej1c2UOdG7SvKwfBUIwWQGfSScDTnrxN3jJY9eGXVxSBGiU9Auh9K8nXyqXv
zqHMmTSa9DM5UlMPyQVWElxNidwF71mY3eAYUXx+IIeSSEfpOsxh4D12D7qEu/VbRGS2NtSL339P
lxLH87Weqpc/om53xkKwuaDihyFgxKptlV/nIst5qT0N3WihAzY/Fu5FI41uIVFkdxBv1VjkLQgL
5kMY+tgUpjdff3u1UuwG15nT1BcHvmJYrfiFC6BDWoLmBZpx2Y5WKFW369C0BQ8zdoa/5e3mT4vV
1XMFoH9hy+2MPrqNLpu5q9+x4JWqtqsVy05SiI2QblPI0g+Wv4B3QlfoRYDuMOz1erxixe17Pgyb
vZDUc0w3WQRSorzDvqDC5/hulFavUWrybQFmW/I6RQPlWkErcKwmSpY5reiWWaMBR1LYbO0lqgiD
K4rTRGOf2pkJ9i/FEkoTHHkyc7kq/G4AAeP5trLqeHS8gssryd6BjJtBYYbBU7RIZwrDUCZ03e0P
NUAR1B1wTkozhMK1WYaLossvI4MiV4SvFAJ82ndGK+sUCduwQ+MqwSZzMwCpwygC4XZQyoFRRm22
CVHYpe+V//RK67UMLlYZCJCD3bOmwOwAUTzimwajbsLYlpprbsKo12M4kXtrTpE59ItxZqVXP/n4
JwH6tr+AIjAJNNaKVcy1v51ZFsPuSdyskqRAB2/H6Hs5jEJ0Pr11pX8F6iBZGDNiuQ4q61d+FRJF
gVA0KSimnDPiznQAudFRHImQz8HCCNzspRAxrwI6qa390pcPOqIC71wnR7AcMC9IH+4kphubD3qn
WhQc0siV7SMzLdYtpQKh0hDBln2ywAw8dWK0lgKyx/DT4Vg7pAng7sAyXUtkhJywVy6cIwetehcv
BxtKRG11ZRdRCirqx0gLvWVBk7bD6fLE2T+QKMDtoPsflIYfOprQI8/ow9gV8k/vaZ5Y6mIHFx7R
+pNGAs9F/6nq9nBNnir+zeNzrli2d1ubBVe/qs/rT4+e0RgxuEIbSdqEFrUlQYU8FCqV9NBzLB2K
8ySCfdrCTDmBEiYIe+fafbMAtKJx9tKWpMkreRelLnZ02po5kCPo0czYQXdCmcUaZv3yIiKRFMSN
x9Lzl0oSKr64jcD1TscOhlEouRurVfSD3cV49qHBOrQEp/cyOyIyut+VeYPoN7ORjlwvSkBhS+0Y
9++sl0vIa6pkqG8AxWseoF6UVkRXBW4Y6JFXM4ynDHrGVG+/Ly063Fd3vjXxXRL+FRbK39oVaoWY
CfnVBZFl2zX7e1ycK+ZZcMD7xSMXNHUI7cBSAEH3P6iwc8/RkYyPpd1cpvzxZG89O1uhbJV5KfIh
Zp3TbV9SZNQJHNpLMPoq2nljzEdib72czZeG6lVKHwtgHLbsmfgYASjB0jyr7LtIXrzXqQUsITEx
3F06O9ARQZ91HfRa7oyibW5gPNCc2oRQ0OsKrJFjERQA0NoIKJxO4TbwAllbGRmkLhAKdDcYDlB/
aM76ClOXIT+mIG5PPhze8Nf8SZOJio6pY8o7bAQyKaNhvPaB4VrlST06c8v2jJR7PysbkUXKAD4j
jmxC7aO5ZHcQliln/Ozz5U1HKrHlZTAL41moDR0EsT33LHpBCO7flFQt8G8WNZauRG5Kl89hMX4E
j7yfc2xCP5NI40Tl/qSC2THeH+PhjE/LKJyaGrKsIVQfaI054faEGYR1yTFg0SwoHZ09tBQrtEor
g8zU1l97e13+76HoPjBzNR3gsp1qTdfSnWrsVPaWiaA0M5N/UniknUjXMzn3Rqn2sgeFF3u+SbS4
QL+tQeKw2SpNY8ZsfPebY+RN1qQbjIai5s3PgwZmgiaFAtjJpa9Ujws3Bnytj9dKR6Qwwwz6iVbd
zrii5FU7Lii8EncZB+bkPCgUxBIwCIC9UkWXPPT9padwcfcpEJCZVvbR0hlGvc7PRZHLRm70veze
QhDKKsDva3clvSDEBp0k6yZ8I6OJ/Z4JZrrl04lJJp3/BaZWMZIXUjyM+/zOvXR08W4gbtsMkJE0
J6gyzQuEhT1o/Vm09rw8fceFwOJg6tb+OcnQ+bTLnrxg2VoQ/X5AjpvHu7wlDJ3M5B0KTLkIKaHP
GEDgEbNq31fjMCEaQ54kX10Mie9ORIqkOd/dDrpAgIb9Tx+A1DkoD7dt3rzqq0usvpCV5Uls1CjT
cW3GBCI14izJB6fEMXXPGdKP5X9xFdMnCoFJ9itBALL9FvsGXrSdF+Qrnvnn7fr8rd9bOgVO02nv
KPZk7yokpaOvRF/Lkv9OmwCYaln4ogmguZYgsOrfFqDoOCEkTPHtYqeIYqCEQoO3DFfMY7i5twVB
FbobFOeGBg/QMJH+OHDWRRcLvM2Yg/LhTPOaJAJ04MrqcAgIUFlAytT2bhxqMsUK18kCvdyrB2Q9
kQ04jqtU3BJeJeSrgdSWRytGt6mBzuj109lUnW7S9ixBZy+CX/Jb/EyZJ5HGhBSb0m7aNSKhItht
sf/GznQRWxO9uK8NvzcDAxCpLn3G5zXMJr4yG3eUSU/bLcNctBo5Qi/qZF66nzrNaDQMpYiOIefI
BR4uBGhZ0rJaBSFewBxrMtktIyOpnoG0R8hr0u6tX8jfpYvnwGFd6kJ9HlkMmY6JvwKl7kYgGQEJ
9vZq1EDWTeSmjDIEGIKwdx51qDHFUqqI83mLmyCFPr9iti19jtzBpra1VGaw265rG+ueEtgvECPZ
uY8R7xo/iBFJPL/YO7m2LpHgpNdxbuC0aCDf5oMRUIiO8Oah4pc2Se9TFie1bjt3EnAC/Ppv3sTP
bT+9/PbsPL8QS373NYLIqVM2o5ZBzAUinD858R8WFi5+PNjconrVdRgZ6avYJSGuFB/XbXcWUErg
S/9VaGa43OT9tfR27j+Pj5ROJqqpcr6hxwsaM9AiDi5QiD5zR5NfSGeix117zwaSZTUTZszCYOAN
7Zz7naPIqbpOqzkkfp0nphRMllTBN3CdG3+VU9byUhEhgvEyp1EEzjhU6iQEx7aKd8ST3B6hjdwD
Ro+5Sv4q4DH8ErFpaPygOONCEky+p59wKe+XDSmuhN81v8dsg2qO5TaprcyDPetwuGQux9xvh06F
ZV10V5Gcu2wGC8XnHX9iwSKQoScNAhWoCMLKDsGedKmoqF3udFr9xPVrsRNxhsa/ZukcLhd/qwUm
Lh0X70lohSpI6H54lBZBFmYOim11mnTovTiy/S+/cSq/1TOXWARs8ZqgindRQorCbgEFP5pvpqMY
5HefXiYKAPwuABENSArWjofSHqw8DvNvpf8+M2EfJZYccfhGhrgOCFrtiw0cSUYVo8DToeCYLzML
zMqS0lBg5L3bUdV4MEg7VqzsjLFxsX02BNhQTTg4obzn1I5CUFvtCSpviY4b3xLslMI8K/Zf71K3
VATFiHtJgmU6n3rQXjPwVHpzRF8xmbF3IswfQNPW+kGrF0HloXlFj0uPZHQB9R0OEGan5cOQXxVf
3A3ZaQdcWQu8wCLyE33HSiUfm5qKTmkerCEQJPQl9Jgj65AzoUGuH5UIa9pPsFM3i9ZqXY6vtSbi
L+WckHbyYALZ6BRMHglapZIYffftAfd/DtMy/Xf/TJfPl8o6TrtmfSibdUvjtPdXkHbQnPrlDjr5
ub/iKPDYjxHXBqyewUqzwU+V4yixUwdWuVBm/I2r5uaz8bO1lrkU85z2dbwIGBI33qe/x4ol3SJu
CbwAq6UQIDUywmu2Pht7A7kIUWZX6Rvz+Ra5oILmLaKiL/+4V9lZf6hkestXY30kHNcFAe2ADQ5n
+tGvJgrcS+bRZ1E05MI+jdZbd/n3kKRlPGAQAbtXCXpfSaF6oXuHaZghqCRiYiN7pggccwDGi5Jf
QxwzFKNe2jraUH6wyu9ziv5XgudF2fDxkuW+TnZrO+bJ12pn8qn5gBcQCFbWqRaC/RKldSaCQEPl
4BRqSOI1odw1XdtkGEjSL4Hug/hYysEs+PaxKGgxmYOjy77CVXTWYAr4Xxj5GjVh1fc6j9xCEQYQ
bYCn4afTEj68t8cz+qdaYyOpg2I2MywE2a5pBWNCp68uyxgN9K/c00DQw7f6f2Xa59G+MW3DcgQX
9Gregxwv0OHlZsSBsmYBOCwdxqzufAK/2wuMaYz/ra9xnEufslNeJdd0UMqPxngCgGta8O+uAEMv
3NcXjX4aWCMBjfzy160lrI9cvnr1pP1SuEBEGOfs5H10Sg63EQ9ajr4q4Boi7NCBZVmTdtFYjzAC
QfYvbDyTOFeihi5/ZXubzaedSjrMF5hiTmWmXJ1Tf/EkqMn4CaO3mnDVsxgig5u6ABEhpxD3HjIB
/FJlxqTqtu6QBYVN4SQvW3ztcZFjQIXysWFM/P6jgIR/rO+NOZvnfUj2tb8pQ2XflzFg0uQXVAcR
r00u06JXgXepUcCw874PX3dFt/v8VOI7fh0bpL3hfSxha39HeczuXUFe55Rvy8MhsrFlLm3MkDV9
cN6TyCRAPDiURx468b73vx6pV8zdEQyYk49vsiYkLdsnPv6+BNzkY+xa95+aO+iF38a+5/c4Q/+8
4NApASg73S3n3c+6aXatC4gNWoBOTAUtNnQWROUoHuoU9xafbp306R1J8JkwzUuaWyyYUysI7Qrv
PuPaPSoZyg20vkUJgyNrkDEvFu2LVOf4JSb2uEr+Zl9yg5siugPPkg+uD8jvIVS+t0qkqcAR4wGt
QmTBb5AfqmWOhaLCJbChr9Jk54OJgys3OTeW5GD3EmtLX+GEwW81rRAwEgpDRZi6HEqXzottAG++
IZEcwkdimN55RtujEE66bvjnEH+mLje2qVn5qSb6F++hNN6ART40lY4GJtP4W1K12zXMGMhojQ85
yPZPWphe3eAl1wh8eeARm2LfXBiVY9fb+ZOW6MFPcLZs+QIHHj7DtL2bl+eS4ndbH/QFEUL9bJzb
HROGosBcJsX9kLUNHlpZz7IjpMIwNmC0Y7uf3lM41C3f2XeUiQV9kXH/ezh0gSYYCk5RlNkZBm+W
xKh2HnY3qVBSDTVsUkiC1ox1LxhC0bkm1fOvVcaqhC8IWCOO6tgaonHuoCP4yCmOzDKkO6SaH2j7
FW4THTQ+N+3YO1+IzXGJmEk9P5IKPh8edGoPxUNQ7WRMie/uO7g6RRV0iAnu0nR/a8Um11HSFXqf
v8NKsNOtSy/wawTfqTZ1gQNU0ztEbTJIRl+sRAvRcNee5yCjCzchO2LF3ykpTAHt1mxazkc7IPQ3
IA4BpmB5M8h6cZZY+LIF5xNm7xs+hJ2pRVzxY+DDN3uY5mN+yuArj56qUFx51f1GnV3LPcd+jlWs
O/fPCZuwRdDc8gzGYIbveGGa0Di0chIVtn4ybavBYC2yGTZ0Bxxg0oVxc6K4Yls0Df7ICHzFWqQH
eVW0ukfWJDSutoUIb1uaHlhYf7v/WE1Gg5lkRpDyByLmTGS5fWvfcMW6T8ZsI7Z+mbur1CkYp0Q0
vcJGgVy+zZiy53N0JspVCCBfnDfSB0llNR995bU/AtoklVKQD0zDGDwbiJD64ufLeF6ZRirmy5e2
N5/dZFnrHcpz2IlY3f7QY3rUfgX80ZL32C1HLjdpYBXXAKMFrgzceKp+xayK/lOcRuDRt/6sqM5w
Sh/C1T+ZJiqLHhweW/mjCoKVUtnnUllmcfGO4p1usG0KBZFEI94lEiC2zzAAVSK11uD21KCQGcER
rLEbA4MBmjYWYTCQRjCveO2ACBLgThmfHr47yWlAz3xNm92zUosyWZK60P1FbvYRKpRFgmtY0mAv
eeRXWpPu9XqpRfRg704CllGz+RXinIKxm2y9nO8b/phUkka8HrrBFPPBawa6CfeHXk0pIxR80j6p
MXM5kgi6NVJsqbpSmf1I5+7gulVJiO3KFmgQ1fC5hMPBDC6oVToFjDtRzwOpVnsRcvGf1DsRD6UT
b2Y4RsSRsEXhkdiD5cWUeC9OwolPgyh9yoy/36fpzXs2XLZSq7abH0ZgEkgRMubaQFchn7wQ4SgD
9sMMYLmhOfj02m/i/doRl5XS9urO2t5VBKXddnC7hLpKpbhTdAM8G9l0/XoDBcvtqOd58SO6rGvU
PIndcOQPvQG6GGLYbmi/0kBalkTZx5DUt1yKzoUFuLINpKbIPdasRSM+sU2NIQhTYgVKwx6PV/Cb
97kji/OAAP9n42eTwZmWJYozy6dvvyhNXJ3PbXYCg4Q5q1nG1b2Wi5EdRu1D1vNQhLBqcYCatXNB
SO56kPQgQwAuyMD4FaD1/gsLE4Uo5rWC3KN+yXyDyDDPCXigGyHhM+pUkP8yHjOB1ttpYAp279zW
CiJyTxv8A9/clnMvqpxpL9F6OeYWF27tIbIxwfAoYRQ6XtnS9cLXG5sepxPytXOtHruzSq1Rg9TW
t+1/Ph1gaPHwg2zEydwvP/u/3bpWrVq8PrXTzF+k/qpiwtqdmwwB4Wjs3YTlDGDezM3mpIC+x8vZ
QrkExQGiueqJT63fxpJczLJFq//15h8dEmL3SVG2PrACl6nS64zwDROrfYrjY7StKADCXZJNgap9
QD8885pyM9LrW8kqppaEsDRwk4dmj5hP5EivjAZj4ZUnDE9Qq91vj3lgG/92urAUi2Ag5b/aJGkh
DgmbPo8XgxLUWXyOUQlAQjJAv7PcXBfcnrGi1kbNaROwoYZkW/xka09r3GN/W+Vta+itBbTyRRl7
6M2Ws0CNxuULURDPQ6y0TJwxGBwP41KqX58P16oNODecNfwCVvkukosXvq7eV4Kg6GywlLYqXiZq
T0+kvnXgybF5MxUioPVKwv8ORPvftduIg+gpVomCJMXvBGlQalL5ulGUESRIANX02LCDK39GQNkW
JsBjD4CDAtlZU9Ya0y/vhhOeKkHT6w7IExyQaERmxR5xxQwPnTe0+Qk57fTsGfoHbSNoTcNSPHZG
MrVs4Gr7gvnlHdvA/UwQTlXUzySu5DJgZI3mGKQQ4k6wuSjd0fxLjUPUl2Shyug0hgxK4HodlCiy
Oenuk8mu0LoDMxHcOcoq0qby2W9lSuiQT1XIXbKIGvQZvOWuoyglA9ML3/LtrmFNhpsKXqUGNW3z
caIATlWHA6XCHZ74QGPhIfx/B3PryLk+rUJQ9t59xW6kr8xz2xppkxRlYMLbRpC0ren6D87jZY5n
IvG+rltxQwNpla3Vz5bFbb8QGtr3ZhXVExBWBJAcHCewopaw5lZ9WfAOkUNyDHf6Yn4PDKz9lzTH
qiuH/K3rOUafOVx8jR55R/cMpRTsWbSfj5UHRUw/C1q8KBLcS0nOHeJYfDtNSwhhwzQD5bv3ZWhA
lmKJo9hpM3p+93ZmuVG/a0Ih9eBA22QV24UX9dY8GNqBd4XHR0pblv7oYogkJFx+Utp6uY18DNqc
bu+Kh9Kt8K6nqy+qzmPdApQn7/cYEvgXIcH5RdraOJaExfVGokkrWPCH02Kbof06vr8/kd4VOTAb
x/n/r/aI+DMN1JMW7NlC2M5wjeYL2eF5u289Om8BthvQswU7q7m9QAbLE2YIiftjadaDYLhaPM2h
gtEoG35pcEDCIyyxrVM0qms83ngYaVffmtE6lpDm2eB9m2pZGTb/PCul7hKB000M2PAET68CG21F
O0No8XfUXEiOyuopxZt6kE/NQxICuCW9JxR7RRCahxYLt6zg1zkte2onshW6FV9KDNQvCBBmYnYf
L7z30RSfe9uRobU6N1OGbmK63pObgQnbDC5i/2XMvfdG1sMdhmnIXoAAqLwdR2VSg47EHJTCX8Ns
OdRQQuxg2VFyQWQbc9Bmp6kafdIxh3g0o++F3xbloSNMh+ydGswKb6Qrv8AVAIN1gsZdncZB6nkd
iSeSvXd7IXChL73ugg2M5zeZJNMQLjtlDkz54UcaWcvPchUi6J7saKnIoMoH/N8Vcqbcp719HvfH
VHvMs4Zb9BPjX8HrQiV5uimKNfZj5XsWAXgqVpflcCsj/daAVpk23uJKGHW0eMYz0fKvKe1QR3c0
2O8eKkPJI3nnIeHLxPnhS4A8DWOGOmoI0nZdPm8pQ28ArVcsjAHx+L5dN3tgQj37bRTbv40CVojX
ShK+hKUSxKmf1voSXAh3OVdbkXQQLUOHER3l/bCZj8YFhUkvPXlT4FIeL2oFpHt+ZPIshmskIl/A
9uCxuilripZnAFGjBBNXu+uQA/ShGWe8o43m4JBagyiZZQXfy3leZGoaABksXyPKd75kaRDqvYTD
Pqyos/WJp5jLmeij35d9f1lQQ/KzG5d0UI/+0btPH/f+MBQWGXddFw0gKtiAAG0YVRi8dyQ6H+fR
drVq/dCMdwbDd194cHYHxeMnr8mJ7CK1tmZNq01Wm08yzkT1b89vkLXUumSjcEiH3sFUWnpv1/pa
FdqgznRJWVLQorZ3KMFs31PWqhpR5H58oCjxmnmS5gL/Q8eKVxJrK48m9I8LDoaftxWs9PcJ7MK2
dHD4laSdUGstxMpBuNlhWVkfJP4b75fvIyT8lfZOVegq8ImEW9lwQXnLzUd8U8xHmhdE40f0xMiD
wJxz94NrOhtdTEKTlYB6EH2sG4SFrA+2WGMBzxe24ieBQNOC7j7IGtKgCrv3TC975qFHQYcFE6pN
CdrHcVZrPGZPV6wM6ReEULrSK5Ikmj7cyW4Z4xBjDLsON6kiA9oiI5dzgdnEqpuz+jYDIGxW4VmP
tv9dSb0ZMWhzD6DD/dxxZpPk8px6FOKJkCRC291AHPX1vNvfUYPIZI6k3tuf1LerPIRBADwI3eTb
sA1/anB6mQEODJaNW02/LCdxlOJx1E0ptN+wPwt+1ws0FkYIcx/PgCjOkzJDQ2iEVew4U/dMrsDX
cYx4//0xa81J6wajLIsQAlqwOpRItRWLtpRd1i6szIiopw55dqQHPmvX6D4svQU223qKQHwk2sdx
x7gLFn7CSdo1fwBbnEvZI8AcgwCqgLXJQxdLIVyCtmph1gTOlnzDXb2xLygHJSGwOrAE0lM8NpU4
e3Kg9m8inlD0F539tsAPPl7yca0ltTUAliMLq53O3k/nbOQFplJE4kQSEQshWxzZeFOxolKkGpru
pSpAEETZnK2qHRFe95brxD8WEWQ/abHulCjG/AakJ/fAuU78fLaeRG3F0GPb/z8Yz/BYbiArqw+Z
GVYiMkkE+uDBecRKj0G+EY+F+Iy9tpz625vv8dGeF/eTbGLRGUS0octtfqfogjPeKIn89VdgMtae
2gDyVWRfCp3wriq0N5b5mo+tqDoSMl5bUnSVNib3YdBF8/llFg+fsOxspBHjx9q1r8qdxjXITfo1
FiDbg2P6ouNQcUKL8C7z7KNwhgvj3OjpYdbeUvOGcbBv5EgEy9iR7vcz1aGnmqWi2/U2vUJ5t2hZ
iRFBYQ7wpMVWajeuu9pUax3B7YSo06zgAKmVvnr8xAwEnr+IFnZ1FRiJ6WQ57DwRE7kr6/Oxxvhp
gE3Cy6SQsZBzLKgr2aXGaZ9HfBWlndthi4eCOvgEcBzK1FxIktpVrciX96LQlEZ+Khw/zpCC0cSf
WLgU8nYe5KRnKUFlCk+JAuNOO/jLlom2fxH61PoLJs9/cO39dhAdsUZQmIs44FRoaVroLIyDxdRB
GEX2gVJ24ntfE9zPs4bmo/r92N4EQZRnUUZEAhO4X8TR1bbfQRGoytCK9NRjFsp3w5/phyPN2hgi
6JkizQM6jDy2KzyfO/aKW6Kz6uIcYzCiVrgSadPbHD/GhnNw6dUErcqnH+dBfJeXZFwioXoI/Yuv
gBHCPRVKlMIgIoUb2t329ynBtWoafpJmBzAUkzNJVIhiEmbavgOcz2GucWn0mJ/lzQVdF9jUBJVq
qqF134ZMa67BRf/P7A+t3jKUOchSdpLMfYqGg/W3ry440lI3W4JO0BCvhYZTvs/S5CTtoGwdM459
tRMyUJwhGzmvwPmcs7NHj6ptjCwOXrco8KRa3OPOZuvibwmNHa+Bydr7zk19Wix7j9mSoJaGLTne
Jk5eQ01o0PYIKtIVOK+IP1A7r+tj6Djm4sSOzN7l/vg0tfePyUy/YuTKyJO+1QCEg45fq3DcPTQg
NMaehNhwMG2iSIK5lYwX/AXVNnRqmrrs9xmX2GB5uMLc2yGcwm+cJq+Q8Ycmn1UgFg74Lj7HiV38
xEpHrdYoYSfg83Xx+ifOAEwFYRPiDGXEUrWsuDBECwUhuNarE0Mqmu2TEFByB7eetbscpGUJzYWU
CvL50M0WMtv+st1G7qkMFwSWo98Oao9IQfHUwwTech4bM5yUAoog9Bo4so3qyRLzkGla7BQsfXZo
1jXokvzFohvwWRMo9ShSLuEM4SOteiMN+P6kU35Q5/t8N3j6HGgCmlgJptzKO/UyIcqEISRP8AGR
/BUJ/EMcgJTrtEG3AmEljwbWL/yY43sdo6IbMclf4RmuPQzcZjhguNfYpoYHnNlRzz0alF8FA746
hG5K97wvWKrc2opYUdsR20cNGcOfsTNsgAYsJzlhOIftjzyDsAe80+q+BV9FW1PDhqfIv7GC/V93
pdgjWbnoxkwp9S8N3EokGDjfHd9gW4uDOtMT5S9Km2xy4K6xpkpeDvfGC7wy3mEujLJHsB1W4mPU
76CHF6MpqRNuhBTMN7uoYLnSfhj4j1iwj1nhxnWy+AaMq2fgFM/diWQZw4UKagi+nSIhVZ1sVouh
CdC8SAgxHyoY8nJn46USN4AKP4W6Hmhd+JGNNyReTNjFNEpLKZE6OFZ7Mrwh8tYS3k72Hs2wxnAl
urejsJ4DDyAEKVTz/T2YC67gtpnQeMyawC4ndwod4xlRfBymYlzG0cCd09LlcTt0v8muEAvz3GXl
jUOodE8tn7mtDKMS4SnDHyePOH4dEjDvbsntMvg8h5CG05uMSBJWbsYBYHKYTvgFutwh+J8pD2ar
GMrbzVR/awNZUoo+Z6YqW0N3S7PxiHHoqzQnuk6RlujKqJkkpyBd2rxr7Mz8K53m08JuA0QCSWLh
5rtDFv6/dYALVXV2jld/pSIr4BJ8TMGLxG2Zf6HxROxGqi7s384LFTUHptqsPl268KNpfU4s7yas
99o9oHwszcnBza0s24biP1fYm4pZ0A34pFYSXUmDyIKfXUbzLpBeWAt62fLxWayhjPkd9BZ+bv+j
7Iz0IB3KmKdP1ABC/ktRjap+KCXNDw1pEElF+QXWm0EWmwJTWzkLyLEqr/KT6uHDeGEGgvQIlKL9
kFT4dOBNwAjLQRkzVyfGHLtfrMoOaphjZIL6tykFmv2xiz6EU0Y2p1g/r+PeLkEbvj6zPdTVjMEK
j1a6rMzlm1DuBx7DMH4m5pE10QM5T06d9xQsZL48vmLDMODeodh/ugzviggPciQaD9TKY7fQnrFR
wuC6uvIfYy1LleaQ0ZdTB6o88Y3ExWicVbkcCLZ+R3v7FJ6KLHHdzpmETxXAFJG4EgmyJu4mZb0x
EBtBTt+54Zjhc7t9CXQQVeemEas1U1mtQLZWVaRG/SB8Fufc3kp6EkoIJgahGGUZEW2YK0ZwszrL
JaXuF0PjJ2TXaEGUuYgLUBjyR2yWliUTWmKHLNwMZeE+E5YfcsuKEoqebt0DY+hsxPu37Q+uBOqJ
qkTcDCKl0mFDQjHq/oS+z92uRQ5uSGdeji9amLQyJMMVI9XvFyvWEFaThlaOXJX1mk52ReiDy1O3
kzrxS8oaY5KHpg8U6v/EShuYs3v1c30Nf82Sxfa2gw7S49/zlxxebLb8OsYFJwtVmnUjc98DsYL5
0GW+PXEW2uCFE5olL81krNTtpcASLCfydLq9CZ1mTLI9zPtRS2sJsiWB2aiQ5y5lCufzHpfRyJuU
PyBu0gvtSxSTX3ellK98XWwjaqYQoR4dTO9fCIkW57/2Zk+TCfm48QYqt7TFtF5uJXZh1QdWfArL
gx95AA8aIRC0y1nhRpT+Wv9F+T0sU/ImwaiDUxvOlOzy9oNWqdzWaEkL2LyvWkV8SuuZj6bmX2bs
OM/jb/vmOyFInih9uGsYpuxQe6kDfJvW9V6Ul9glAEhdBOOm8w6EW6LLBQXhOuelMLqqy0clN6mv
k44evMPcI59c+N+RFSR7lzyvlwnJrBSRh3HpLnywTBjUYSUfo3yKrtsnq1QynYmmQXPy+JAdmND0
+YrHmLJrjyvQKuGVLAVsF9Yjd0Y7lAD2G3KKFMjtG3qiGt+KLUygwAod6nuAj0DTRgS4n+XDV/yN
YBHueLECsJRYIqKKpMU0B9etnEVi0//fBs6BW8xwio1bWc7aYqOOdv3/bZPP43/feoQ9o5a3FuJS
S9FNouW4M1fg+NbtIhESwMTyivebuDg8Piqz1uHGRqGt6EOGtTNER+vc6JFUOzxfLiVnpyLcWyxz
GCr7wNBsixMTxq/oTgHKcXD38kqA06VQNr1qIoFPXlprGhBQWHx95RNfXOJn1aOatMeGUnvzqSEu
FPK/LZky+VQUNxBC2coBzu7HHY4nVV8EjScpQokjDgHegkuALU+Og6udf4tmHIAQL8GmB9amWmhq
y70JfW365lGt4OSrK5tIVdSKxa/qdyoSn3Fc91f8qLXQlAxm6rCX/q5Kov310/gG35qIJErGiNT6
HyKK9fOVZWMNsfoiANdadzDfyJkuOpEb0968ESnXaNBbzdZEV/nsWtC+/YjtoGFd9seVopEO7RxI
zvMHS4vwccpVMuXMYsL6LTokdGL2+CiHVzVX4u0DNGwfa1o7pepWiovPA5VNmqgVyfYw6eeixFoq
wJNzN9HBZUPE/UtvYlZ5IfzFIvaviior0B+tTWVstN0wlY8yQm9m6e6tqq43zeLz+EJr+Q4y3JdY
8l2U8VD1uoggRD2Yd3+tL/uV8QnoGEMub3+hexC6g3vNb2UJLESDUZ2IwfCUdAHU1OSzybGQ4elL
pc5qPHIZH8jZbo4da4Xf7Qx3frYAd67iFnPlIpZ9ACNxcVdD7KtT9O4EUUVowXPYw1/SGUWUTiZ6
+kdqy21leD15DVWCZYtG6nt0/8ofp04evxBlS6Eux8tGO4vftvPQ7wGHXpAG6SqLwBtiHD/noDmQ
j6jvW/2rDiXvc6rxzPALTE+wQ5zu3lgSZhYpC3WevmbMAncJp1L3XacJrfRHJVrRpRwpHzI1o7uX
4DF/3yUstxI5YsgVDMyQIaSDUEHlTl0z/LJog/803Z7EIBYh05EIVTa1NEkvgLsPWnejZ3T9kV9G
vXjC9tEpGSrnmel9jOxVORG6Byu0+zo5Tkiz7VntVAYWVE3/5S2fLk7Y0WMC6gc+GUhX3WkWm94C
7ow5mDLUHYdEPZncatg3UggJy17K2wnXcVRllanQSs3zQWcxmZmJ0ZkPh2jC2TtT97aW4etb0Xyb
EY4YOqmh/huf63UITST+Bt2DjsUMlJbeH6Ja6s2n7i77+flK/PpiLicE1z+PmZ2/Sh01ILScCNQW
uDpUCkRFCm5wYk8puSs3sFlsa08BpI1xdISlPDhUgtv69I/6
`protect end_protected
